//#### BEGIN MODULE DEFINITION FOR :AFIFO36_INTERNAL ###
module AFIFO36_INTERNAL (ALMOSTEMPTY, ALMOSTFULL, DBITERR, DO, DOP, ECCPARITY, EMPTY, FULL, RDCOUNT, RDERR, SBITERR, WRCOUNT, WRERR,
			DI, DIP, RDCLK, RDEN, RDRCLK, RST, WRCLK, WREN) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [63:0] DI ;
input [7:0] DIP ;
input RDCLK ;
input RDEN ;
input RDRCLK ;
input RST ;
input WRCLK ;
input WREN ;
output ALMOSTEMPTY ;
output ALMOSTFULL ;
output DBITERR ;
output [63:0] DO ;
output [7:0] DOP ;
output [7:0] ECCPARITY ;
output EMPTY ;
output FULL ;
output [12:0] RDCOUNT ;
output RDERR ;
output SBITERR ;
output [12:0] WRCOUNT ;
output WRERR ;
parameter DATA_WIDTH = 4;
parameter DO_REG = 1;
parameter EN_SYN = "FALSE";
parameter FIRST_WORD_FALL_THROUGH = "FALSE";
parameter ALMOST_EMPTY_OFFSET = 13'h0080;
parameter ALMOST_FULL_OFFSET = 13'h0080;
parameter EN_ECC_WRITE = "FALSE";
parameter EN_ECC_READ = "FALSE";
parameter SIM_MODE = "SAFE";
parameter FIFO_SIZE = 36;
endmodule
//#### END MODULE DEFINITION FOR: AFIFO36_INTERNAL ####

//#### BEGIN MODULE DEFINITION FOR :AND2 ###
module AND2 (O, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND2 ####

//#### BEGIN MODULE DEFINITION FOR :AND2B1 ###
module AND2B1 (O, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND2B1 ####

//#### BEGIN MODULE DEFINITION FOR :AND2B1L ###
module AND2B1L (O,  DI, SRI) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input SRI ;
input DI ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND2B1L ####

//#### BEGIN MODULE DEFINITION FOR :AND2B2 ###
module AND2B2 (O, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND2B2 ####

//#### BEGIN MODULE DEFINITION FOR :AND3 ###
module AND3 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND3 ####

//#### BEGIN MODULE DEFINITION FOR :AND3B1 ###
module AND3B1 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND3B1 ####

//#### BEGIN MODULE DEFINITION FOR :AND3B2 ###
module AND3B2 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND3B2 ####

//#### BEGIN MODULE DEFINITION FOR :AND3B3 ###
module AND3B3 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND3B3 ####

//#### BEGIN MODULE DEFINITION FOR :AND4 ###
module AND4 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND4 ####

//#### BEGIN MODULE DEFINITION FOR :AND4B1 ###
module AND4B1 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND4B1 ####

//#### BEGIN MODULE DEFINITION FOR :AND4B2 ###
module AND4B2 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND4B2 ####

//#### BEGIN MODULE DEFINITION FOR :AND4B3 ###
module AND4B3 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND4B3 ####

//#### BEGIN MODULE DEFINITION FOR :AND4B4 ###
module AND4B4 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND4B4 ####

//#### BEGIN MODULE DEFINITION FOR :AND5 ###
module AND5 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND5 ####

//#### BEGIN MODULE DEFINITION FOR :AND5B1 ###
module AND5B1 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND5B1 ####

//#### BEGIN MODULE DEFINITION FOR :AND5B2 ###
module AND5B2 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND5B2 ####

//#### BEGIN MODULE DEFINITION FOR :AND5B3 ###
module AND5B3 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND5B3 ####

//#### BEGIN MODULE DEFINITION FOR :AND5B4 ###
module AND5B4 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND5B4 ####

//#### BEGIN MODULE DEFINITION FOR :AND5B5 ###
module AND5B5 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: AND5B5 ####

//#### BEGIN MODULE DEFINITION FOR :ARAMB36_INTERNAL ###
module ARAMB36_INTERNAL (CASCADEOUTLATA, CASCADEOUTLATB, CASCADEOUTREGA, CASCADEOUTREGB, DBITERR, DOA, DOB, DOPA, DOPB, ECCPARITY, SBITERR, 
			 ADDRA, ADDRB, CASCADEINLATA, CASCADEINLATB, CASCADEINREGA, CASCADEINREGB, CLKA, CLKB, DIA, DIB, DIPA, DIPB, ENA, ENB, GSR, REGCEA, REGCEB, REGCLKA, REGCLKB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input ENA ;
input CLKA ;
input REGCLKA ;
input SSRA ;
input CASCADEINLATA ;
input CASCADEINREGA ;
input REGCEA ;
input ENB ;
input CLKB ;
input REGCLKB ;
input SSRB ;
input CASCADEINLATB ;
input CASCADEINREGB ;
input REGCEB ;
input GSR ;
input [15:0] ADDRA ;
input [15:0] ADDRB ;
input [63:0] DIA ;
input [63:0] DIB ;
input [3:0] DIPA ;
input [7:0] DIPB ;
input [7:0] WEA ;
input [7:0] WEB ;
output CASCADEOUTLATA ;
output CASCADEOUTREGA ;
output CASCADEOUTLATB ;
output CASCADEOUTREGB ;
output SBITERR ;
output DBITERR ;
output [63:0] DOA ;
output [31:0] DOB ;
output [7:0] DOPA ;
output [3:0] DOPB ;
output [7:0] ECCPARITY ;
parameter DOA_REG = 0;
parameter DOB_REG = 0;
parameter EN_ECC_READ = "FALSE";
parameter EN_ECC_SCRUB = "FALSE";
parameter EN_ECC_WRITE = "FALSE";
parameter INIT_A = 72'h0;
parameter INIT_B = 72'h0;
parameter RAM_EXTENSION_A = "NONE";
parameter RAM_EXTENSION_B = "NONE";
parameter READ_WIDTH_A = 0;
parameter READ_WIDTH_B = 0;
parameter SETUP_ALL = 1000;
parameter SETUP_READ_FIRST = 3000;
parameter SIM_COLLISION_CHECK = "ALL";
parameter SRVAL_A = 72'h0;
parameter SRVAL_B = 72'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter WRITE_WIDTH_A = 0;
parameter WRITE_WIDTH_B = 0;
parameter INIT_FILE = "NONE";
parameter SIM_MODE = "SAFE";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_40 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_41 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_42 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_43 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_44 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_45 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_46 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_47 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_48 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_49 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_50 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_51 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_52 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_53 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_54 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_55 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_56 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_57 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_58 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_59 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_60 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_61 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_62 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_63 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_64 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_65 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_66 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_67 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_68 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_69 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_70 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_71 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_72 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_73 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_74 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_75 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_76 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_77 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_78 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_79 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter BRAM_MODE = "TRUE_DUAL_PORT";
parameter BRAM_SIZE = 36;
endmodule
//#### END MODULE DEFINITION FOR: ARAMB36_INTERNAL ####

//#### BEGIN MODULE DEFINITION FOR :AUTOBUF ###
module AUTOBUF (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
parameter BUFFER_TYPE = "AUTO";
endmodule
//#### END MODULE DEFINITION FOR: AUTOBUF ####

//#### BEGIN MODULE DEFINITION FOR :BSCANE2 ###
module BSCANE2 (
  CAPTURE,
  DRCK,
  RESET,
  RUNTEST,
  SEL,
  SHIFT,
  TCK,
  TDI,
  TMS,
  UPDATE,

  TDO
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input TDO ;
output CAPTURE ;
output DRCK ;
output RESET ;
output RUNTEST ;
output SEL ;
output SHIFT ;
output TCK ;
output TDI ;
output TMS ;
output UPDATE ;
parameter DISABLE_JTAG = "FALSE";
parameter JTAG_CHAIN = 1;
endmodule
//#### END MODULE DEFINITION FOR: BSCANE2 ####

//#### BEGIN MODULE DEFINITION FOR :BSCAN_FPGACORE ###
module BSCAN_FPGACORE (CAPTURE, DRCK1, DRCK2, RESET, SEL1, SEL2, SHIFT, TDI, UPDATE, TDO1, TDO2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input TDO1 ;
input TDO2 ;
output CAPTURE ;
output DRCK1 ;
output DRCK2 ;
output RESET ;
output SEL1 ;
output SEL2 ;
output SHIFT ;
output TDI ;
output UPDATE ;
endmodule
//#### END MODULE DEFINITION FOR: BSCAN_FPGACORE ####

//#### BEGIN MODULE DEFINITION FOR :BSCAN_SPARTAN3 ###
module BSCAN_SPARTAN3 (CAPTURE, DRCK1, DRCK2, RESET, SEL1, SEL2, SHIFT, TDI, UPDATE, TDO1, TDO2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input TDO1 ;
input TDO2 ;
output CAPTURE ;
output DRCK1 ;
output DRCK2 ;
output RESET ;
output SEL1 ;
output SEL2 ;
output SHIFT ;
output TDI ;
output UPDATE ;
endmodule
//#### END MODULE DEFINITION FOR: BSCAN_SPARTAN3 ####

//#### BEGIN MODULE DEFINITION FOR :BSCAN_SPARTAN3A ###
module BSCAN_SPARTAN3A (CAPTURE, DRCK1, DRCK2, RESET, SEL1, SEL2, SHIFT, TCK, TDI, TMS, UPDATE, TDO1, TDO2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input TDO1 ;
input TDO2 ;
output CAPTURE ;
output DRCK1 ;
output DRCK2 ;
output RESET ;
output SEL1 ;
output SEL2 ;
output SHIFT ;
output TCK ;
output TDI ;
output TMS ;
output UPDATE ;
endmodule
//#### END MODULE DEFINITION FOR: BSCAN_SPARTAN3A ####

//#### BEGIN MODULE DEFINITION FOR :BSCAN_SPARTAN6 ###
module BSCAN_SPARTAN6 (CAPTURE, DRCK, RESET, RUNTEST, SEL, SHIFT, TCK, TDI, TMS, UPDATE, TDO) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input TDO ;
output CAPTURE ;
output DRCK ;
output RESET ;
output RUNTEST ;
output SEL ;
output SHIFT ;
output TCK ;
output TDI ;
output TMS ;
output UPDATE ;
parameter JTAG_CHAIN = 1;
endmodule
//#### END MODULE DEFINITION FOR: BSCAN_SPARTAN6 ####

//#### BEGIN MODULE DEFINITION FOR :BSCAN_VIRTEX4 ###
module BSCAN_VIRTEX4 (CAPTURE, DRCK, RESET, SEL, SHIFT, TDI, UPDATE, TDO) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input TDO ;
output CAPTURE ;
output DRCK ;
output RESET ;
output SEL ;
output SHIFT ;
output TDI ;
output UPDATE ;
parameter JTAG_CHAIN = 1;
endmodule
//#### END MODULE DEFINITION FOR: BSCAN_VIRTEX4 ####

//#### BEGIN MODULE DEFINITION FOR :BSCAN_VIRTEX5 ###
module BSCAN_VIRTEX5 (CAPTURE, DRCK, RESET, SEL, SHIFT, TDI, UPDATE, TDO) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input TDO ;
output CAPTURE ;
output DRCK ;
output RESET ;
output SEL ;
output SHIFT ;
output TDI ;
output UPDATE ;
parameter JTAG_CHAIN = 1;
endmodule
//#### END MODULE DEFINITION FOR: BSCAN_VIRTEX5 ####

//#### BEGIN MODULE DEFINITION FOR :BSCAN_VIRTEX6 ###
module BSCAN_VIRTEX6 (
  CAPTURE,
  DRCK,
  RESET,
  RUNTEST,
  SEL,
  SHIFT,
  TCK,
  TDI,
  TMS,
  UPDATE,
  TDO
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input TDO ;
output CAPTURE ;
output DRCK ;
output RESET ;
output RUNTEST ;
output SEL ;
output SHIFT ;
output TCK ;
output TDI ;
output TMS ;
output UPDATE ;
parameter DISABLE_JTAG = "FALSE";
parameter JTAG_CHAIN = 1;
endmodule
//#### END MODULE DEFINITION FOR: BSCAN_VIRTEX6 ####

//#### BEGIN MODULE DEFINITION FOR :BUF ###
module BUF (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: BUF ####

//#### BEGIN MODULE DEFINITION FOR :BUFCF ###
module BUFCF (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: BUFCF ####

//#### BEGIN MODULE DEFINITION FOR :BUFE ###
module BUFE (O, E, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input E ;
input I ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: BUFE ####

//#### BEGIN MODULE DEFINITION FOR :BUFG ###
module BUFG (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: BUFG ####

//#### BEGIN MODULE DEFINITION FOR :BUFGCE ###
module BUFGCE (O, CE, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CE ;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: BUFGCE ####

//#### BEGIN MODULE DEFINITION FOR :BUFGCE_1 ###
module BUFGCE_1 (O, CE, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CE ;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: BUFGCE_1 ####

//#### BEGIN MODULE DEFINITION FOR :BUFGCTRL ###
module BUFGCTRL (O, CE0, CE1, I0, I1, IGNORE0, IGNORE1, S0, S1) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CE0 ;
input CE1 ;
input I0 ;
input I1 ;
input IGNORE0 ;
input IGNORE1 ;
input S0 ;
input S1 ;
output O ;
parameter INIT_OUT = 0;
parameter PRESELECT_I0 = "FALSE";
parameter PRESELECT_I1 = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: BUFGCTRL ####

//#### BEGIN MODULE DEFINITION FOR :BUFGDLL ###
module BUFGDLL (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
parameter DUTY_CYCLE_CORRECTION = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: BUFGDLL ####

//#### BEGIN MODULE DEFINITION FOR :BUFGMUX ###
module BUFGMUX (O, I0, I1, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input S ;
output O ;
parameter CLK_SEL_TYPE = "SYNC";
endmodule
//#### END MODULE DEFINITION FOR: BUFGMUX ####

//#### BEGIN MODULE DEFINITION FOR :BUFGMUX_1 ###
module BUFGMUX_1 (O, I0, I1, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input S ;
output O ;
parameter CLK_SEL_TYPE = "SYNC";
endmodule
//#### END MODULE DEFINITION FOR: BUFGMUX_1 ####

//#### BEGIN MODULE DEFINITION FOR :BUFGMUX_CTRL ###
module BUFGMUX_CTRL (O, I0, I1, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input S ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: BUFGMUX_CTRL ####

//#### BEGIN MODULE DEFINITION FOR :BUFGMUX_VIRTEX4 ###
module BUFGMUX_VIRTEX4 (O, I0, I1, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input S ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: BUFGMUX_VIRTEX4 ####

//#### BEGIN MODULE DEFINITION FOR :BUFGP ###
module BUFGP (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: BUFGP ####

//#### BEGIN MODULE DEFINITION FOR :BUFG_LB ###
module BUFG_LB (
  CLKOUT,

  CLKIN
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKIN ;
output CLKOUT ;
endmodule
//#### END MODULE DEFINITION FOR: BUFG_LB ####

//#### BEGIN MODULE DEFINITION FOR :BUFH ###
module BUFH (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: BUFH ####

//#### BEGIN MODULE DEFINITION FOR :BUFHCE ###
module BUFHCE (O, CE, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CE ;
input I ;
output O ;
parameter CE_TYPE = "SYNC";
parameter INIT_OUT = 0;
endmodule
//#### END MODULE DEFINITION FOR: BUFHCE ####

//#### BEGIN MODULE DEFINITION FOR :BUFIO ###
module BUFIO (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: BUFIO ####

//#### BEGIN MODULE DEFINITION FOR :BUFIO2 ###
module BUFIO2 (DIVCLK, IOCLK, SERDESSTROBE, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output DIVCLK ;
output IOCLK ;
output SERDESSTROBE ;
parameter DIVIDE_BYPASS = "TRUE";
parameter DIVIDE = 1;
parameter I_INVERT = "FALSE";
parameter USE_DOUBLER = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: BUFIO2 ####

//#### BEGIN MODULE DEFINITION FOR :BUFIO2FB ###
module BUFIO2FB (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
parameter DIVIDE_BYPASS = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: BUFIO2FB ####

//#### BEGIN MODULE DEFINITION FOR :BUFIO2_2CLK ###
module BUFIO2_2CLK (DIVCLK, IOCLK, SERDESSTROBE, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output DIVCLK ;
output IOCLK ;
output SERDESSTROBE ;
parameter DIVIDE = 2;
endmodule
//#### END MODULE DEFINITION FOR: BUFIO2_2CLK ####

//#### BEGIN MODULE DEFINITION FOR :BUFIODQS ###
module BUFIODQS (O, DQSMASK, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input DQSMASK ;
input I ;
output O ;
parameter DQSMASK_ENABLE = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: BUFIODQS ####

//#### BEGIN MODULE DEFINITION FOR :BUFMR ###
module BUFMR (
  O,

  I
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: BUFMR ####

//#### BEGIN MODULE DEFINITION FOR :BUFMRCE ###
module BUFMRCE (
  O,

  CE,
  I
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CE ;
input I ;
output O ;
parameter CE_TYPE = "SYNC";
parameter INIT_OUT = 0;
endmodule
//#### END MODULE DEFINITION FOR: BUFMRCE ####

//#### BEGIN MODULE DEFINITION FOR :BUFPLL ###
module BUFPLL (IOCLK, LOCK, SERDESSTROBE, GCLK, LOCKED, PLLIN) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input GCLK ;
input LOCKED ;
input PLLIN ;
output IOCLK ;
output LOCK ;
output SERDESSTROBE ;
parameter DIVIDE = 1;
parameter ENABLE_SYNC = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: BUFPLL ####

//#### BEGIN MODULE DEFINITION FOR :BUFPLL_MCB ###
module BUFPLL_MCB (
  IOCLK0,
  IOCLK1,
  LOCK,
  SERDESSTROBE0,
  SERDESSTROBE1,

  GCLK,
  LOCKED,
  PLLIN0,
  PLLIN1
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input GCLK ;
input LOCKED ;
input PLLIN0 ;
input PLLIN1 ;
output IOCLK0 ;
output IOCLK1 ;
output LOCK ;
output SERDESSTROBE0 ;
output SERDESSTROBE1 ;
parameter DIVIDE = 2;
parameter LOCK_SRC = "LOCK_TO_0";
endmodule
//#### END MODULE DEFINITION FOR: BUFPLL_MCB ####

//#### BEGIN MODULE DEFINITION FOR :BUFR ###
module BUFR (O, CE, CLR, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CE ;
input CLR ;
input I ;
output O ;
parameter BUFR_DIVIDE = "BYPASS";
parameter SIM_DEVICE = "VIRTEX4";
endmodule
//#### END MODULE DEFINITION FOR: BUFR ####

//#### BEGIN MODULE DEFINITION FOR :BUFT ###
module BUFT (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: BUFT ####

//#### BEGIN MODULE DEFINITION FOR :CAPTUREE2 ###
module CAPTUREE2 (
  CAP,
  CLK
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CAP ;
input CLK ;
parameter ONESHOT = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: CAPTUREE2 ####

//#### BEGIN MODULE DEFINITION FOR :CAPTURE_FPGACORE ###
module CAPTURE_FPGACORE (CAP, CLK) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CAP ;
input CLK ;
parameter ONESHOT = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: CAPTURE_FPGACORE ####

//#### BEGIN MODULE DEFINITION FOR :CAPTURE_SPARTAN3 ###
module CAPTURE_SPARTAN3 (CAP, CLK) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CAP ;
input CLK ;
parameter ONESHOT = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: CAPTURE_SPARTAN3 ####

//#### BEGIN MODULE DEFINITION FOR :CAPTURE_SPARTAN3A ###
module CAPTURE_SPARTAN3A (CAP, CLK) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CAP ;
input CLK ;
parameter ONESHOT = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: CAPTURE_SPARTAN3A ####

//#### BEGIN MODULE DEFINITION FOR :CAPTURE_VIRTEX4 ###
module CAPTURE_VIRTEX4 (CAP, CLK) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CAP ;
input CLK ;
parameter ONESHOT = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: CAPTURE_VIRTEX4 ####

//#### BEGIN MODULE DEFINITION FOR :CAPTURE_VIRTEX5 ###
module CAPTURE_VIRTEX5 (
	CAP,
	CLK
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CAP ;
input CLK ;
parameter ONESHOT = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: CAPTURE_VIRTEX5 ####

//#### BEGIN MODULE DEFINITION FOR :CAPTURE_VIRTEX6 ###
module CAPTURE_VIRTEX6 (
  CAP,
  CLK
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CAP ;
input CLK ;
parameter ONESHOT = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: CAPTURE_VIRTEX6 ####

//#### BEGIN MODULE DEFINITION FOR :CARRY4 ###
module CARRY4 (CO, O, CI, CYINIT, DI, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CI ;
input CYINIT ;
input [3:0] DI ;
input [3:0] S ;
output [3:0] CO ;
output [3:0] O ;
endmodule
//#### END MODULE DEFINITION FOR: CARRY4 ####

//#### BEGIN MODULE DEFINITION FOR :CFGLUT5 ###
module CFGLUT5 (CDO, O5, O6, CDI, CE, CLK, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I4 ;
input I3 ;
input I2 ;
input I1 ;
input I0 ;
input CDI ;
input CE ;
input CLK ;
output CDO ;
output O5 ;
output O6 ;
parameter INIT = 32'h00000000;
endmodule
//#### END MODULE DEFINITION FOR: CFGLUT5 ####

//#### BEGIN MODULE DEFINITION FOR :CLKDLL ###
module CLKDLL (
	CLK0, CLK180, CLK270, CLK2X, CLK90, CLKDV, LOCKED, 
	CLKFB, CLKIN, RST) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKFB ;
input CLKIN ;
input RST ;
output CLK0 ;
output CLK180 ;
output CLK270 ;
output CLK2X ;
output CLK90 ;
output CLKDV ;
output LOCKED ;
parameter CLKDV_DIVIDE = 2.0;
parameter DUTY_CYCLE_CORRECTION = "TRUE";
parameter FACTORY_JF = 16'hC080;
parameter STARTUP_WAIT = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: CLKDLL ####

//#### BEGIN MODULE DEFINITION FOR :CLKDLLE ###
module CLKDLLE (
	CLK0, CLK180, CLK270, CLK2X, CLK2X180, CLK90, CLKDV, LOCKED, 
	CLKFB, CLKIN, RST) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKFB ;
input CLKIN ;
input RST ;
output CLK0 ;
output CLK180 ;
output CLK270 ;
output CLK2X ;
output CLK2X180 ;
output CLK90 ;
output CLKDV ;
output LOCKED ;
parameter CLKDV_DIVIDE = 2.0;
parameter DUTY_CYCLE_CORRECTION = "TRUE";
parameter FACTORY_JF = 16'hC080;
parameter STARTUP_WAIT = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: CLKDLLE ####

//#### BEGIN MODULE DEFINITION FOR :CLKDLLHF ###
module CLKDLLHF (
	CLK0, CLK180, CLKDV, LOCKED, 
	CLKFB, CLKIN, RST) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKFB ;
input CLKIN ;
input RST ;
output CLK0 ;
output CLK180 ;
output CLKDV ;
output LOCKED ;
parameter CLKDV_DIVIDE = 2.0;
parameter DUTY_CYCLE_CORRECTION = "TRUE";
parameter FACTORY_JF = 16'hFFF0;
parameter STARTUP_WAIT = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: CLKDLLHF ####

//#### BEGIN MODULE DEFINITION FOR :CONFIG ###
module CONFIG () /* synthesis syn_black_box  syn_lib_cell=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: CONFIG ####

//#### BEGIN MODULE DEFINITION FOR :CRC32 ###
module CRC32 (CRCOUT,
	      CRCCLK,
	      CRCDATAVALID,
	      CRCDATAWIDTH,
	      CRCIN,
	      CRCRESET
	      ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CRCCLK ;
input CRCDATAVALID ;
input [2:0] 	 CRCDATAWIDTH ;
input [31:0]  CRCIN ;
input CRCRESET ;
output [31:0] CRCOUT ;
parameter CRC_INIT = 32'hFFFFFFFF;
endmodule
//#### END MODULE DEFINITION FOR: CRC32 ####

//#### BEGIN MODULE DEFINITION FOR :CRC64 ###
module CRC64 (
	      CRCOUT,
	      CRCCLK,
	      CRCDATAVALID,
	      CRCDATAWIDTH,
	      CRCIN,
	      CRCRESET
	      ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CRCCLK ;
input CRCDATAVALID ;
input [2:0] 	 CRCDATAWIDTH ;
input [63:0]  CRCIN ;
input CRCRESET ;
output [31:0] CRCOUT ;
parameter CRC_INIT = 32'hFFFFFFFF;
endmodule
//#### END MODULE DEFINITION FOR: CRC64 ####

//#### BEGIN MODULE DEFINITION FOR :DCIRESET ###
module DCIRESET (LOCKED, RST) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input RST ;
output LOCKED ;
endmodule
//#### END MODULE DEFINITION FOR: DCIRESET ####

//#### BEGIN MODULE DEFINITION FOR :DCM ###
module DCM (
	CLK0, CLK180, CLK270, CLK2X, CLK2X180, CLK90,
	CLKDV, CLKFX, CLKFX180, LOCKED, PSDONE, STATUS,
	CLKFB, CLKIN, DSSEN, PSCLK, PSEN, PSINCDEC, RST) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKFB ;
input CLKIN ;
input DSSEN ;
input PSCLK ;
input PSEN ;
input PSINCDEC ;
input RST ;
output CLK0 ;
output CLK180 ;
output CLK270 ;
output CLK2X ;
output CLK2X180 ;
output CLK90 ;
output CLKDV ;
output CLKFX ;
output CLKFX180 ;
output LOCKED ;
output PSDONE ;
output [7:0] STATUS ;
parameter CLKDV_DIVIDE = 2.0;
parameter CLKFX_DIVIDE = 1;
parameter CLKFX_MULTIPLY = 4;
parameter CLKIN_DIVIDE_BY_2 = "FALSE";
parameter CLKIN_PERIOD = 10.0;
parameter CLKOUT_PHASE_SHIFT = "NONE";
parameter CLK_FEEDBACK = "1X";
parameter DESKEW_ADJUST = "SYSTEM_SYNCHRONOUS";
parameter DFS_FREQUENCY_MODE = "LOW";
parameter DLL_FREQUENCY_MODE = "LOW";
parameter DSS_MODE = "NONE";
parameter DUTY_CYCLE_CORRECTION = "TRUE";
parameter FACTORY_JF = 16'hC080;
parameter PHASE_SHIFT = 0;
parameter SIM_MODE = "SAFE";
parameter STARTUP_WAIT = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: DCM ####

//#### BEGIN MODULE DEFINITION FOR :DCM_ADV ###
module DCM_ADV (
        CLK0,
        CLK180,
        CLK270,
        CLK2X,
        CLK2X180,
        CLK90,
        CLKDV,
        CLKFX,
        CLKFX180,
        DO,
        DRDY,
        LOCKED,
        PSDONE,
        CLKFB,
        CLKIN,
        DADDR,
        DCLK,
        DEN,
        DI,
        DWE,
        PSCLK,
        PSEN,
        PSINCDEC,
        RST
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKFB ;
input CLKIN ;
input DCLK ;
input DEN ;
input DWE ;
input PSCLK ;
input PSEN ;
input PSINCDEC ;
input RST ;
input [15:0] DI ;
input [6:0] DADDR ;
output CLK0 ;
output CLK180 ;
output CLK270 ;
output CLK2X180 ;
output CLK2X ;
output CLK90 ;
output CLKDV ;
output CLKFX180 ;
output CLKFX ;
output DRDY ;
output LOCKED ;
output PSDONE ;
output [15:0] DO ;
parameter CLKDV_DIVIDE = 2.0;
parameter CLKFX_DIVIDE = 1;
parameter CLKFX_MULTIPLY = 4;
parameter CLKIN_DIVIDE_BY_2 = "FALSE";
parameter CLKIN_PERIOD = 10.0;
parameter CLKOUT_PHASE_SHIFT = "NONE";
parameter CLK_FEEDBACK = "1X";
parameter DCM_AUTOCALIBRATION = "TRUE";
parameter DCM_PERFORMANCE_MODE = "MAX_SPEED";
parameter DESKEW_ADJUST = "SYSTEM_SYNCHRONOUS";
parameter DFS_FREQUENCY_MODE = "LOW";
parameter DLL_FREQUENCY_MODE = "LOW";
parameter DUTY_CYCLE_CORRECTION = "TRUE";
parameter FACTORY_JF = 16'hF0F0;
parameter PHASE_SHIFT = 0;
parameter SIM_DEVICE ="VIRTEX4";
parameter STARTUP_WAIT = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: DCM_ADV ####

//#### BEGIN MODULE DEFINITION FOR :DCM_BASE ###
module DCM_BASE (
	CLK0,
	CLK180,
	CLK270,
	CLK2X,
	CLK2X180,
	CLK90,
	CLKDV,
	CLKFX,
	CLKFX180,
	LOCKED,
	CLKFB,
	CLKIN,
	RST
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKFB ;
input CLKIN ;
input RST ;
output CLK0 ;
output CLK180 ;
output CLK270 ;
output CLK2X180 ;
output CLK2X ;
output CLK90 ;
output CLKDV ;
output CLKFX180 ;
output CLKFX ;
output LOCKED ;
parameter CLKDV_DIVIDE = 2.0;
parameter CLKFX_DIVIDE = 1;
parameter CLKFX_MULTIPLY = 4;
parameter CLKIN_DIVIDE_BY_2 = "FALSE";
parameter CLKIN_PERIOD = 10.0;
parameter CLKOUT_PHASE_SHIFT = "NONE";
parameter CLK_FEEDBACK = "1X";
parameter DCM_AUTOCALIBRATION = "TRUE";
parameter DCM_PERFORMANCE_MODE = "MAX_SPEED";
parameter DESKEW_ADJUST = "SYSTEM_SYNCHRONOUS";
parameter DFS_FREQUENCY_MODE = "LOW";
parameter DLL_FREQUENCY_MODE = "LOW";
parameter DUTY_CYCLE_CORRECTION = "TRUE";
parameter FACTORY_JF = 16'hF0F0;
parameter PHASE_SHIFT = 0;
parameter STARTUP_WAIT = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: DCM_BASE ####

//#### BEGIN MODULE DEFINITION FOR :DCM_CLKGEN ###
module DCM_CLKGEN (
  CLKFX,
  CLKFX180,
  CLKFXDV,
  LOCKED,
  PROGDONE,
  STATUS,
  CLKIN,
  FREEZEDCM,
  PROGCLK,
  PROGDATA,
  PROGEN,
  RST
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKIN ;
input FREEZEDCM ;
input PROGCLK ;
input PROGDATA ;
input PROGEN ;
input RST ;
output CLKFX180 ;
output CLKFX ;
output CLKFXDV ;
output LOCKED ;
output PROGDONE ;
output [2:1] STATUS ;
parameter SPREAD_SPECTRUM = "NONE";
parameter STARTUP_WAIT = "FALSE";
parameter CLKFXDV_DIVIDE = 2;
parameter CLKFX_DIVIDE = 1;
parameter CLKFX_MULTIPLY = 4;
parameter CLKFX_MD_MAX = 0.0;
parameter CLKIN_PERIOD = 0.0;
endmodule
//#### END MODULE DEFINITION FOR: DCM_CLKGEN ####

//#### BEGIN MODULE DEFINITION FOR :DCM_PS ###
module DCM_PS (
	CLK0,
	CLK180,
	CLK270,
	CLK2X,
	CLK2X180,
	CLK90,
	CLKDV,
	CLKFX,
	CLKFX180,
	DO,
	LOCKED,
	PSDONE,
	CLKFB,
	CLKIN,
	PSCLK,
	PSEN,
	PSINCDEC,
	RST
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKFB ;
input CLKIN ;
input PSCLK ;
input PSEN ;
input PSINCDEC ;
input RST ;
output CLK0 ;
output CLK180 ;
output CLK270 ;
output CLK2X180 ;
output CLK2X ;
output CLK90 ;
output CLKDV ;
output CLKFX180 ;
output CLKFX ;
output LOCKED ;
output PSDONE ;
output [15:0] DO ;
parameter CLKDV_DIVIDE = 2.0;
parameter CLKFX_DIVIDE = 1;
parameter CLKFX_MULTIPLY = 4;
parameter CLKIN_DIVIDE_BY_2 = "FALSE";
parameter CLKIN_PERIOD = 10.0;
parameter CLKOUT_PHASE_SHIFT = "NONE";
parameter CLK_FEEDBACK = "1X";
parameter DCM_AUTOCALIBRATION = "TRUE";
parameter DCM_PERFORMANCE_MODE = "MAX_SPEED";
parameter DESKEW_ADJUST = "SYSTEM_SYNCHRONOUS";
parameter DFS_FREQUENCY_MODE = "LOW";
parameter DLL_FREQUENCY_MODE = "LOW";
parameter DUTY_CYCLE_CORRECTION = "TRUE";
parameter FACTORY_JF = 16'hF0F0;
parameter PHASE_SHIFT = 0;
parameter STARTUP_WAIT = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: DCM_PS ####

//#### BEGIN MODULE DEFINITION FOR :DCM_SP ###
module DCM_SP (
	CLK0, CLK180, CLK270, CLK2X, CLK2X180, CLK90,
	CLKDV, CLKFX, CLKFX180, LOCKED, PSDONE, STATUS,
	CLKFB, CLKIN, DSSEN, PSCLK, PSEN, PSINCDEC, RST) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKFB ;
input CLKIN ;
input DSSEN ;
input PSCLK ;
input PSEN ;
input PSINCDEC ;
input RST ;
output CLK0 ;
output CLK180 ;
output CLK270 ;
output CLK2X ;
output CLK2X180 ;
output CLK90 ;
output CLKDV ;
output CLKFX ;
output CLKFX180 ;
output LOCKED ;
output PSDONE ;
output [7:0] STATUS ;
parameter CLKDV_DIVIDE = 2.0;
parameter CLKFX_DIVIDE = 1;
parameter CLKFX_MULTIPLY = 4;
parameter CLKIN_DIVIDE_BY_2 = "FALSE";
parameter CLKIN_PERIOD = 10.0;
parameter CLKOUT_PHASE_SHIFT = "NONE";
parameter CLK_FEEDBACK = "1X";
parameter DESKEW_ADJUST = "SYSTEM_SYNCHRONOUS";
parameter DFS_FREQUENCY_MODE = "LOW";
parameter DLL_FREQUENCY_MODE = "LOW";
parameter DSS_MODE = "NONE";
parameter DUTY_CYCLE_CORRECTION = "TRUE";
parameter FACTORY_JF = 16'hC080;
parameter PHASE_SHIFT = 0;
parameter STARTUP_WAIT = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: DCM_SP ####

//#### BEGIN MODULE DEFINITION FOR :DNA_PORT ###
module DNA_PORT (DOUT, CLK, DIN, READ, SHIFT) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLK ;
input DIN ;
input READ ;
input SHIFT ;
output DOUT ;
parameter SIM_DNA_VALUE = 57'h0;
endmodule
//#### END MODULE DEFINITION FOR: DNA_PORT ####

//#### BEGIN MODULE DEFINITION FOR :DSP48 ###
module DSP48 (BCOUT, P, PCOUT, A, B, BCIN, C, CARRYIN, CARRYINSEL, CEA, CEB, CEC, CECARRYIN, CECINSUB, CECTRL, CEM, CEP, CLK, OPMODE, PCIN, RSTA, RSTB, RSTC, RSTCARRYIN, RSTCTRL, RSTM, RSTP, SUBTRACT)  /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [17:0] A ;
input [17:0] B ;
input [17:0] BCIN ;
input [47:0] C ;
input CARRYIN ;
input [1:0] CARRYINSEL ;
input CEA ;
input CEB ;
input CEC ;
input CECARRYIN ;
input CECINSUB ;
input CECTRL ;
input CEM ;
input CEP ;
input CLK ;
input [6:0] OPMODE ;
input [47:0] PCIN ;
input RSTA ;
input RSTB ;
input RSTC ;
input RSTCARRYIN ;
input RSTCTRL ;
input RSTM ;
input RSTP ;
input SUBTRACT ;
output [17:0] BCOUT ;
output [47:0] P ;
output [47:0] PCOUT ;
parameter AREG = 1;
parameter BREG = 1;
parameter B_INPUT = "DIRECT";
parameter CARRYINREG = 1;
parameter CARRYINSELREG = 1;
parameter CREG = 1;
parameter LEGACY_MODE = "MULT18X18S";
parameter MREG = 1;
parameter OPMODEREG = 1;
parameter PREG = 1;
parameter SUBTRACTREG = 1;
endmodule
//#### END MODULE DEFINITION FOR: DSP48 ####

//#### BEGIN MODULE DEFINITION FOR :DSP48A ###
module DSP48A (BCOUT, CARRYOUT, P, PCOUT, A, B, C, CARRYIN, CEA, CEB, CEC, CECARRYIN, CED, CEM, CEOPMODE, CEP, CLK, D, OPMODE, PCIN, RSTA, RSTB, RSTC, RSTCARRYIN, RSTD, RSTM, RSTOPMODE, RSTP)  /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [17:0] A ;
input [17:0] B ;
input [47:0] C ;
input CARRYIN ;
input CEA ;
input CEB ;
input CEC ;
input CECARRYIN ;
input CED ;
input CEM ;
input CEOPMODE ;
input CEP ;
input CLK ;
input [17:0] D ;
input [7:0] OPMODE ;
input [47:0] PCIN ;
input RSTA ;
input RSTB ;
input RSTC ;
input RSTCARRYIN ;
input RSTD ;
input RSTM ;
input RSTOPMODE ;
input RSTP ;
output [17:0] BCOUT ;
output CARRYOUT ;
output [47:0] P ;
output [47:0] PCOUT ;
parameter A0REG = 0;
parameter A1REG = 1;
parameter B0REG = 0;
parameter B1REG = 1;
parameter CARRYINREG = 1;
parameter CARRYINSEL = "CARRYIN";
parameter CREG = 1;
parameter DREG = 1;
parameter MREG = 1;
parameter OPMODEREG = 1;
parameter PREG = 1;
parameter RSTTYPE = "SYNC";
endmodule
//#### END MODULE DEFINITION FOR: DSP48A ####

//#### BEGIN MODULE DEFINITION FOR :DSP48A1 ###
module DSP48A1 (BCOUT, CARRYOUT, CARRYOUTF, M, P, PCOUT, A, B, C, CARRYIN, CEA, CEB, CEC, CECARRYIN, CED, CEM, CEOPMODE, CEP, CLK, D, OPMODE, PCIN, RSTA, RSTB, RSTC, RSTCARRYIN, RSTD, RSTM, RSTOPMODE, RSTP)  /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [17:0] A ;
input [17:0] B ;
input [47:0] C ;
input CARRYIN ;
input CEA ;
input CEB ;
input CEC ;
input CECARRYIN ;
input CED ;
input CEM ;
input CEOPMODE ;
input CEP ;
input CLK ;
input [17:0] D ;
input [7:0] OPMODE ;
input [47:0] PCIN ;
input RSTA ;
input RSTB ;
input RSTC ;
input RSTCARRYIN ;
input RSTD ;
input RSTM ;
input RSTOPMODE ;
input RSTP ;
output [17:0] BCOUT ;
output CARRYOUT ;
output CARRYOUTF ;
output [35:0] M ;
output [47:0] P ;
output [47:0] PCOUT ;
parameter A0REG = 0;
parameter A1REG = 1;
parameter B0REG = 0;
parameter B1REG = 1;
parameter CARRYINREG = 1;
parameter CARRYOUTREG = 1;
parameter CARRYINSEL = "OPMODE5";
parameter CREG = 1;
parameter DREG = 1;
parameter MREG = 1;
parameter OPMODEREG = 1;
parameter PREG = 1;
parameter RSTTYPE = "SYNC";
endmodule
//#### END MODULE DEFINITION FOR: DSP48A1 ####

//#### BEGIN MODULE DEFINITION FOR :DSP48E ###
module DSP48E (ACOUT, BCOUT, CARRYCASCOUT, CARRYOUT, MULTSIGNOUT, OVERFLOW, P, PATTERNBDETECT, PATTERNDETECT, PCOUT, UNDERFLOW, A, ACIN, ALUMODE, B, BCIN, C, CARRYCASCIN, CARRYIN, CARRYINSEL, CEA1, CEA2, CEALUMODE, CEB1, CEB2, CEC, CECARRYIN, CECTRL, CEM, CEMULTCARRYIN, CEP, CLK, MULTSIGNIN, OPMODE, PCIN, RSTA, RSTALLCARRYIN, RSTALUMODE, RSTB, RSTC, RSTCTRL, RSTM, RSTP)  /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [29:0] A ;
input [29:0] ACIN ;
input [3:0] ALUMODE ;
input [17:0] B ;
input [17:0] BCIN ;
input [47:0] C ;
input CARRYCASCIN ;
input CARRYIN ;
input [2:0] CARRYINSEL ;
input CEA1 ;
input CEA2 ;
input CEALUMODE ;
input CEB1 ;
input CEB2 ;
input CEC ;
input CECARRYIN ;
input CECTRL ;
input CEM ;
input CEMULTCARRYIN ;
input CEP ;
input CLK ;
input MULTSIGNIN ;
input [6:0] OPMODE ;
input [47:0] PCIN ;
input RSTA ;
input RSTALLCARRYIN ;
input RSTALUMODE ;
input RSTB ;
input RSTC ;
input RSTCTRL ;
input RSTM ;
input RSTP ;
output [29:0] ACOUT ;
output [17:0] BCOUT ;
output CARRYCASCOUT ;
output [3:0] CARRYOUT ;
output MULTSIGNOUT ;
output OVERFLOW ;
output [47:0] P ;
output PATTERNBDETECT ;
output PATTERNDETECT ;
output [47:0] PCOUT ;
output UNDERFLOW ;
parameter SIM_MODE = "SAFE";
parameter ACASCREG = 1;
parameter ALUMODEREG = 1;
parameter AREG = 1;
parameter AUTORESET_PATTERN_DETECT = "FALSE";
parameter AUTORESET_PATTERN_DETECT_OPTINV = "MATCH";
parameter A_INPUT = "DIRECT";
parameter BCASCREG = 1;
parameter BREG = 1;
parameter B_INPUT = "DIRECT";
parameter CARRYINREG = 1;
parameter CARRYINSELREG = 1;
parameter CREG = 1;
parameter MASK =  48'h3FFFFFFFFFFF;
parameter MREG = 1;
parameter MULTCARRYINREG = 1;
parameter OPMODEREG = 1;
parameter PATTERN =  48'h000000000000;
parameter PREG = 1;
parameter SEL_MASK = "MASK";
parameter SEL_PATTERN = "PATTERN";
parameter SEL_ROUNDING_MASK = "SEL_MASK";
parameter USE_MULT = "MULT_S";
parameter USE_PATTERN_DETECT = "NO_PATDET";
parameter USE_SIMD = "ONE48";
endmodule
//#### END MODULE DEFINITION FOR: DSP48E ####

//#### BEGIN MODULE DEFINITION FOR :DSP48E1 ###
module DSP48E1 (ACOUT, BCOUT, CARRYCASCOUT, CARRYOUT, MULTSIGNOUT, OVERFLOW, P, PATTERNBDETECT, PATTERNDETECT, PCOUT, UNDERFLOW, A, ACIN, ALUMODE, B, BCIN, C, CARRYCASCIN, CARRYIN, CARRYINSEL, CEA1, CEA2, CEAD, CEALUMODE, CEB1, CEB2, CEC, CECARRYIN, CECTRL, CED, CEINMODE, CEM, CEP, CLK, D, INMODE, MULTSIGNIN, OPMODE, PCIN, RSTA, RSTALLCARRYIN, RSTALUMODE, RSTB, RSTC, RSTCTRL, RSTD, RSTINMODE, RSTM, RSTP)  /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [29:0] A ;
input [29:0] ACIN ;
input [3:0] ALUMODE ;
input [17:0] B ;
input [17:0] BCIN ;
input [47:0] C ;
input CARRYCASCIN ;
input CARRYIN ;
input [2:0] CARRYINSEL ;
input CEA1 ;
input CEA2 ;
input CEAD ;
input CEALUMODE ;
input CEB1 ;
input CEB2 ;
input CEC ;
input CECARRYIN ;
input CECTRL ;
input CED ;
input CEINMODE ;
input CEM ;
input CEP ;
input CLK ;
input [24:0] D ;
input [4:0] INMODE ;
input MULTSIGNIN ;
input [6:0] OPMODE ;
input [47:0] PCIN ;
input RSTA ;
input RSTALLCARRYIN ;
input RSTALUMODE ;
input RSTB ;
input RSTC ;
input RSTCTRL ;
input RSTD ;
input RSTINMODE ;
input RSTM ;
input RSTP ;
output [29:0] ACOUT ;
output [17:0] BCOUT ;
output CARRYCASCOUT ;
output [3:0] CARRYOUT ;
output MULTSIGNOUT ;
output OVERFLOW ;
output [47:0] P ;
output PATTERNBDETECT ;
output PATTERNDETECT ;
output [47:0] PCOUT ;
output UNDERFLOW ;
parameter ACASCREG = 1;
parameter ADREG = 1;
parameter ALUMODEREG = 1;
parameter AREG = 1;
parameter AUTORESET_PATDET = "NO_RESET";
parameter A_INPUT = "DIRECT";
parameter BCASCREG = 1;
parameter BREG = 1;
parameter B_INPUT = "DIRECT";
parameter CARRYINREG = 1;
parameter CARRYINSELREG = 1;
parameter CREG = 1;
parameter DREG = 1;
parameter INMODEREG = 1;
parameter MASK =  48'h3FFFFFFFFFFF;
parameter MREG = 1;
parameter OPMODEREG = 1;
parameter PATTERN =  48'h000000000000;
parameter PREG = 1;
parameter SEL_MASK = "MASK";
parameter SEL_PATTERN = "PATTERN";
parameter USE_DPORT = "FALSE";
parameter USE_MULT = "MULTIPLY";
parameter USE_PATTERN_DETECT = "NO_PATDET";
parameter USE_SIMD = "ONE48";
endmodule
//#### END MODULE DEFINITION FOR: DSP48E1 ####

//#### BEGIN MODULE DEFINITION FOR :DSP48E2 ###
module DSP48E2 (ACOUT, BCOUT, CARRYCASCOUT, CARRYOUT, MULTSIGNOUT, OVERFLOW, P, PATTERNBDETECT, PATTERNDETECT, PCOUT, UNDERFLOW, XORTREE, A, ACIN, ALUMODE, B, BCIN, C, CARRYCASCIN, CARRYIN, CARRYINSEL, CEA1, CEA2, CEAD, CEALUMODE, CEB1, CEB2, CEC, CECARRYIN, CECTRL, CED, CEINMODE, CEM, CEP, CLK, D, INMODE, MULTSIGNIN, OPMODE, PCIN, RSTA, RSTALLCARRYIN, RSTALUMODE, RSTB, RSTC, RSTCTRL, RSTD, RSTINMODE, RSTM, RSTP)  /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [29:0] A ;
input [29:0] ACIN ;
input [3:0] ALUMODE ;
input [17:0] B ;
input [17:0] BCIN ;
input [47:0] C ;
input CARRYCASCIN ;
input CARRYIN ;
input [2:0] CARRYINSEL ;
input CEA1 ;
input CEA2 ;
input CEAD ;
input CEALUMODE ;
input CEB1 ;
input CEB2 ;
input CEC ;
input CECARRYIN ;
input CECTRL ;
input CED ;
input CEINMODE ;
input CEM ;
input CEP ;
input CLK ;
input [26:0] D ;
input [4:0] INMODE ;
input MULTSIGNIN ;
input [8:0] OPMODE ;
input [47:0] PCIN ;
input RSTA ;
input RSTALLCARRYIN ;
input RSTALUMODE ;
input RSTB ;
input RSTC ;
input RSTCTRL ;
input RSTD ;
input RSTINMODE ;
input RSTM ;
input RSTP ;
output [29:0] ACOUT ;
output [17:0] BCOUT ;
output CARRYCASCOUT ;
output [3:0] CARRYOUT ;
output MULTSIGNOUT ;
output OVERFLOW ;
output [47:0] P ;
output PATTERNBDETECT ;
output PATTERNDETECT ;
output [47:0] PCOUT ;
output UNDERFLOW ;
output [7:0] XORTREE;
parameter ACASCREG = 1;
parameter ADREG = 1;
parameter ALUMODEREG = 1;
parameter AREG = 1;
parameter AUTORESET_PATDET = "NO_RESET";
parameter A_INPUT = "DIRECT";
parameter BCASCREG = 1;
parameter BREG = 1;
parameter B_INPUT = "DIRECT";
parameter CARRYINREG = 1;
parameter CARRYINSELREG = 1;
parameter CREG = 1;
parameter DREG = 1;
parameter INMODEREG = 1;
parameter MASK =  48'h3FFFFFFFFFFF;
parameter MREG = 1;
parameter OPMODEREG = 1;
parameter PATTERN =  48'h000000000000;
parameter PREG = 1;
parameter SEL_MASK = "MASK";
parameter SEL_PATTERN = "PATTERN";
parameter AMULTSEL = "A";
parameter USE_MULT = "MULTIPLY";
parameter USE_PATTERN_DETECT = "NO_PATDET";
parameter USE_SIMD = "ONE48";
parameter RND =  48'h000000000000;
parameter XOR_SIMD = "ONE96";
parameter PREADDINSEL = 0;
parameter BMULTSEL = "B";
endmodule
//#### END MODULE DEFINITION FOR: DSP48E2 ####

//#### BEGIN MODULE DEFINITION FOR :EFUSE_USR ###
module EFUSE_USR (
  EFUSEUSR
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
output [31:0] EFUSEUSR ;
parameter [31:0] SIM_EFUSE_VALUE = 32'h00000000;
endmodule
//#### END MODULE DEFINITION FOR: EFUSE_USR ####

//#### BEGIN MODULE DEFINITION FOR :EMAC ###
module EMAC (
	DCRHOSTDONEIR,
	EMAC0CLIENTANINTERRUPT,
	EMAC0CLIENTRXBADFRAME,
	EMAC0CLIENTRXCLIENTCLKOUT,
	EMAC0CLIENTRXD,
	EMAC0CLIENTRXDVLD,
	EMAC0CLIENTRXDVLDMSW,
	EMAC0CLIENTRXDVREG6,
	EMAC0CLIENTRXFRAMEDROP,
	EMAC0CLIENTRXGOODFRAME,
	EMAC0CLIENTRXSTATS,
	EMAC0CLIENTRXSTATSBYTEVLD,
	EMAC0CLIENTRXSTATSVLD,
	EMAC0CLIENTTXACK,
	EMAC0CLIENTTXCLIENTCLKOUT,
	EMAC0CLIENTTXCOLLISION,
	EMAC0CLIENTTXGMIIMIICLKOUT,
	EMAC0CLIENTTXRETRANSMIT,
	EMAC0CLIENTTXSTATS,
	EMAC0CLIENTTXSTATSBYTEVLD,
	EMAC0CLIENTTXSTATSVLD,
	EMAC0PHYENCOMMAALIGN,
	EMAC0PHYLOOPBACKMSB,
	EMAC0PHYMCLKOUT,
	EMAC0PHYMDOUT,
	EMAC0PHYMDTRI,
	EMAC0PHYMGTRXRESET,
	EMAC0PHYMGTTXRESET,
	EMAC0PHYPOWERDOWN,
	EMAC0PHYSYNCACQSTATUS,
	EMAC0PHYTXCHARDISPMODE,
	EMAC0PHYTXCHARDISPVAL,
	EMAC0PHYTXCHARISK,
	EMAC0PHYTXCLK,
	EMAC0PHYTXD,
	EMAC0PHYTXEN,
	EMAC0PHYTXER,
	EMAC1CLIENTANINTERRUPT,
	EMAC1CLIENTRXBADFRAME,
	EMAC1CLIENTRXCLIENTCLKOUT,
	EMAC1CLIENTRXD,
	EMAC1CLIENTRXDVLD,
	EMAC1CLIENTRXDVLDMSW,
	EMAC1CLIENTRXDVREG6,
	EMAC1CLIENTRXFRAMEDROP,
	EMAC1CLIENTRXGOODFRAME,
	EMAC1CLIENTRXSTATS,
	EMAC1CLIENTRXSTATSBYTEVLD,
	EMAC1CLIENTRXSTATSVLD,
	EMAC1CLIENTTXACK,
	EMAC1CLIENTTXCLIENTCLKOUT,
	EMAC1CLIENTTXCOLLISION,
	EMAC1CLIENTTXGMIIMIICLKOUT,
	EMAC1CLIENTTXRETRANSMIT,
	EMAC1CLIENTTXSTATS,
	EMAC1CLIENTTXSTATSBYTEVLD,
	EMAC1CLIENTTXSTATSVLD,
	EMAC1PHYENCOMMAALIGN,
	EMAC1PHYLOOPBACKMSB,
	EMAC1PHYMCLKOUT,
	EMAC1PHYMDOUT,
	EMAC1PHYMDTRI,
	EMAC1PHYMGTRXRESET,
	EMAC1PHYMGTTXRESET,
	EMAC1PHYPOWERDOWN,
	EMAC1PHYSYNCACQSTATUS,
	EMAC1PHYTXCHARDISPMODE,
	EMAC1PHYTXCHARDISPVAL,
	EMAC1PHYTXCHARISK,
	EMAC1PHYTXCLK,
	EMAC1PHYTXD,
	EMAC1PHYTXEN,
	EMAC1PHYTXER,
	EMACDCRACK,
	EMACDCRDBUS,
	HOSTMIIMRDY,
	HOSTRDDATA,
	CLIENTEMAC0DCMLOCKED,
	CLIENTEMAC0PAUSEREQ,
	CLIENTEMAC0PAUSEVAL,
	CLIENTEMAC0RXCLIENTCLKIN,
	CLIENTEMAC0TXCLIENTCLKIN,
	CLIENTEMAC0TXD,
	CLIENTEMAC0TXDVLD,
	CLIENTEMAC0TXDVLDMSW,
	CLIENTEMAC0TXFIRSTBYTE,
	CLIENTEMAC0TXGMIIMIICLKIN,
	CLIENTEMAC0TXIFGDELAY,
	CLIENTEMAC0TXUNDERRUN,
	CLIENTEMAC1DCMLOCKED,
	CLIENTEMAC1PAUSEREQ,
	CLIENTEMAC1PAUSEVAL,
	CLIENTEMAC1RXCLIENTCLKIN,
	CLIENTEMAC1TXCLIENTCLKIN,
	CLIENTEMAC1TXD,
	CLIENTEMAC1TXDVLD,
	CLIENTEMAC1TXDVLDMSW,
	CLIENTEMAC1TXFIRSTBYTE,
	CLIENTEMAC1TXGMIIMIICLKIN,
	CLIENTEMAC1TXIFGDELAY,
	CLIENTEMAC1TXUNDERRUN,
	DCREMACABUS,
	DCREMACCLK,
	DCREMACDBUS,
	DCREMACENABLE,
	DCREMACREAD,
	DCREMACWRITE,
	HOSTADDR,
	HOSTCLK,
	HOSTEMAC1SEL,
	HOSTMIIMSEL,
	HOSTOPCODE,
	HOSTREQ,
	HOSTWRDATA,
	PHYEMAC0COL,
	PHYEMAC0CRS,
	PHYEMAC0GTXCLK,
	PHYEMAC0MCLKIN,
	PHYEMAC0MDIN,
	PHYEMAC0MIITXCLK,
	PHYEMAC0PHYAD,
	PHYEMAC0RXBUFERR,
	PHYEMAC0RXBUFSTATUS,
	PHYEMAC0RXCHARISCOMMA,
	PHYEMAC0RXCHARISK,
	PHYEMAC0RXCHECKINGCRC,
	PHYEMAC0RXCLK,
	PHYEMAC0RXCLKCORCNT,
	PHYEMAC0RXCOMMADET,
	PHYEMAC0RXD,
	PHYEMAC0RXDISPERR,
	PHYEMAC0RXDV,
	PHYEMAC0RXER,
	PHYEMAC0RXLOSSOFSYNC,
	PHYEMAC0RXNOTINTABLE,
	PHYEMAC0RXRUNDISP,
	PHYEMAC0SIGNALDET,
	PHYEMAC0TXBUFERR,
	PHYEMAC1COL,
	PHYEMAC1CRS,
	PHYEMAC1GTXCLK,
	PHYEMAC1MCLKIN,
	PHYEMAC1MDIN,
	PHYEMAC1MIITXCLK,
	PHYEMAC1PHYAD,
	PHYEMAC1RXBUFERR,
	PHYEMAC1RXBUFSTATUS,
	PHYEMAC1RXCHARISCOMMA,
	PHYEMAC1RXCHARISK,
	PHYEMAC1RXCHECKINGCRC,
	PHYEMAC1RXCLK,
	PHYEMAC1RXCLKCORCNT,
	PHYEMAC1RXCOMMADET,
	PHYEMAC1RXD,
	PHYEMAC1RXDISPERR,
	PHYEMAC1RXDV,
	PHYEMAC1RXER,
	PHYEMAC1RXLOSSOFSYNC,
	PHYEMAC1RXNOTINTABLE,
	PHYEMAC1RXRUNDISP,
	PHYEMAC1SIGNALDET,
	PHYEMAC1TXBUFERR,
	RESET,
	TIEEMAC0CONFIGVEC,
	TIEEMAC0UNICASTADDR,
	TIEEMAC1CONFIGVEC,
	TIEEMAC1UNICASTADDR
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLIENTEMAC0DCMLOCKED ;
input CLIENTEMAC0PAUSEREQ ;
input CLIENTEMAC0RXCLIENTCLKIN ;
input CLIENTEMAC0TXCLIENTCLKIN ;
input CLIENTEMAC0TXDVLD ;
input CLIENTEMAC0TXDVLDMSW ;
input CLIENTEMAC0TXFIRSTBYTE ;
input CLIENTEMAC0TXGMIIMIICLKIN ;
input CLIENTEMAC0TXUNDERRUN ;
input CLIENTEMAC1DCMLOCKED ;
input CLIENTEMAC1PAUSEREQ ;
input CLIENTEMAC1RXCLIENTCLKIN ;
input CLIENTEMAC1TXCLIENTCLKIN ;
input CLIENTEMAC1TXDVLD ;
input CLIENTEMAC1TXDVLDMSW ;
input CLIENTEMAC1TXFIRSTBYTE ;
input CLIENTEMAC1TXGMIIMIICLKIN ;
input CLIENTEMAC1TXUNDERRUN ;
input DCREMACCLK ;
input DCREMACENABLE ;
input DCREMACREAD ;
input DCREMACWRITE ;
input HOSTCLK ;
input HOSTEMAC1SEL ;
input HOSTMIIMSEL ;
input HOSTREQ ;
input PHYEMAC0COL ;
input PHYEMAC0CRS ;
input PHYEMAC0GTXCLK ;
input PHYEMAC0MCLKIN ;
input PHYEMAC0MDIN ;
input PHYEMAC0MIITXCLK ;
input PHYEMAC0RXBUFERR ;
input PHYEMAC0RXCHARISCOMMA ;
input PHYEMAC0RXCHARISK ;
input PHYEMAC0RXCHECKINGCRC ;
input PHYEMAC0RXCLK ;
input PHYEMAC0RXCOMMADET ;
input PHYEMAC0RXDISPERR ;
input PHYEMAC0RXDV ;
input PHYEMAC0RXER ;
input PHYEMAC0RXNOTINTABLE ;
input PHYEMAC0RXRUNDISP ;
input PHYEMAC0SIGNALDET ;
input PHYEMAC0TXBUFERR ;
input PHYEMAC1COL ;
input PHYEMAC1CRS ;
input PHYEMAC1GTXCLK ;
input PHYEMAC1MCLKIN ;
input PHYEMAC1MDIN ;
input PHYEMAC1MIITXCLK ;
input PHYEMAC1RXBUFERR ;
input PHYEMAC1RXCHARISCOMMA ;
input PHYEMAC1RXCHARISK ;
input PHYEMAC1RXCHECKINGCRC ;
input PHYEMAC1RXCLK ;
input PHYEMAC1RXCOMMADET ;
input PHYEMAC1RXDISPERR ;
input PHYEMAC1RXDV ;
input PHYEMAC1RXER ;
input PHYEMAC1RXNOTINTABLE ;
input PHYEMAC1RXRUNDISP ;
input PHYEMAC1SIGNALDET ;
input PHYEMAC1TXBUFERR ;
input RESET ;
input [0:31] DCREMACDBUS ;
input [15:0] CLIENTEMAC0PAUSEVAL ;
input [15:0] CLIENTEMAC0TXD ;
input [15:0] CLIENTEMAC1PAUSEVAL ;
input [15:0] CLIENTEMAC1TXD ;
input [1:0] HOSTOPCODE ;
input [1:0] PHYEMAC0RXBUFSTATUS ;
input [1:0] PHYEMAC0RXLOSSOFSYNC ;
input [1:0] PHYEMAC1RXBUFSTATUS ;
input [1:0] PHYEMAC1RXLOSSOFSYNC ;
input [2:0] PHYEMAC0RXCLKCORCNT ;
input [2:0] PHYEMAC1RXCLKCORCNT ;
input [31:0] HOSTWRDATA ;
input [47:0] TIEEMAC0UNICASTADDR ;
input [47:0] TIEEMAC1UNICASTADDR ;
input [4:0] PHYEMAC0PHYAD ;
input [4:0] PHYEMAC1PHYAD ;
input [79:0] TIEEMAC0CONFIGVEC ;
input [79:0] TIEEMAC1CONFIGVEC ;
input [7:0] CLIENTEMAC0TXIFGDELAY ;
input [7:0] CLIENTEMAC1TXIFGDELAY ;
input [7:0] PHYEMAC0RXD ;
input [7:0] PHYEMAC1RXD ;
input [8:9] DCREMACABUS ;
input [9:0] HOSTADDR ;
output DCRHOSTDONEIR ;
output EMAC0CLIENTANINTERRUPT ;
output EMAC0CLIENTRXBADFRAME ;
output EMAC0CLIENTRXCLIENTCLKOUT ;
output EMAC0CLIENTRXDVLD ;
output EMAC0CLIENTRXDVLDMSW ;
output EMAC0CLIENTRXDVREG6 ;
output EMAC0CLIENTRXFRAMEDROP ;
output EMAC0CLIENTRXGOODFRAME ;
output EMAC0CLIENTRXSTATSBYTEVLD ;
output EMAC0CLIENTRXSTATSVLD ;
output EMAC0CLIENTTXACK ;
output EMAC0CLIENTTXCLIENTCLKOUT ;
output EMAC0CLIENTTXCOLLISION ;
output EMAC0CLIENTTXGMIIMIICLKOUT ;
output EMAC0CLIENTTXRETRANSMIT ;
output EMAC0CLIENTTXSTATS ;
output EMAC0CLIENTTXSTATSBYTEVLD ;
output EMAC0CLIENTTXSTATSVLD ;
output EMAC0PHYENCOMMAALIGN ;
output EMAC0PHYLOOPBACKMSB ;
output EMAC0PHYMCLKOUT ;
output EMAC0PHYMDOUT ;
output EMAC0PHYMDTRI ;
output EMAC0PHYMGTRXRESET ;
output EMAC0PHYMGTTXRESET ;
output EMAC0PHYPOWERDOWN ;
output EMAC0PHYSYNCACQSTATUS ;
output EMAC0PHYTXCHARDISPMODE ;
output EMAC0PHYTXCHARDISPVAL ;
output EMAC0PHYTXCHARISK ;
output EMAC0PHYTXCLK ;
output EMAC0PHYTXEN ;
output EMAC0PHYTXER ;
output EMAC1CLIENTANINTERRUPT ;
output EMAC1CLIENTRXBADFRAME ;
output EMAC1CLIENTRXCLIENTCLKOUT ;
output EMAC1CLIENTRXDVLD ;
output EMAC1CLIENTRXDVLDMSW ;
output EMAC1CLIENTRXDVREG6 ;
output EMAC1CLIENTRXFRAMEDROP ;
output EMAC1CLIENTRXGOODFRAME ;
output EMAC1CLIENTRXSTATSBYTEVLD ;
output EMAC1CLIENTRXSTATSVLD ;
output EMAC1CLIENTTXACK ;
output EMAC1CLIENTTXCLIENTCLKOUT ;
output EMAC1CLIENTTXCOLLISION ;
output EMAC1CLIENTTXGMIIMIICLKOUT ;
output EMAC1CLIENTTXRETRANSMIT ;
output EMAC1CLIENTTXSTATS ;
output EMAC1CLIENTTXSTATSBYTEVLD ;
output EMAC1CLIENTTXSTATSVLD ;
output EMAC1PHYENCOMMAALIGN ;
output EMAC1PHYLOOPBACKMSB ;
output EMAC1PHYMCLKOUT ;
output EMAC1PHYMDOUT ;
output EMAC1PHYMDTRI ;
output EMAC1PHYMGTRXRESET ;
output EMAC1PHYMGTTXRESET ;
output EMAC1PHYPOWERDOWN ;
output EMAC1PHYSYNCACQSTATUS ;
output EMAC1PHYTXCHARDISPMODE ;
output EMAC1PHYTXCHARDISPVAL ;
output EMAC1PHYTXCHARISK ;
output EMAC1PHYTXCLK ;
output EMAC1PHYTXEN ;
output EMAC1PHYTXER ;
output EMACDCRACK ;
output HOSTMIIMRDY ;
output [0:31] EMACDCRDBUS ;
output [15:0] EMAC0CLIENTRXD ;
output [15:0] EMAC1CLIENTRXD ;
output [31:0] HOSTRDDATA ;
output [6:0] EMAC0CLIENTRXSTATS ;
output [6:0] EMAC1CLIENTRXSTATS ;
output [7:0] EMAC0PHYTXD ;
output [7:0] EMAC1PHYTXD ;
endmodule
//#### END MODULE DEFINITION FOR: EMAC ####

//#### BEGIN MODULE DEFINITION FOR :FD ###
module FD (Q, C, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input D ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FD ####

//#### BEGIN MODULE DEFINITION FOR :FDC ###
module FDC (Q, C, CLR, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CLR ;
input D ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDC ####

//#### BEGIN MODULE DEFINITION FOR :FDCE ###
module FDCE (Q, C, CE, CLR, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input CLR ;
input D ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDCE ####

//#### BEGIN MODULE DEFINITION FOR :FDCE_1 ###
module FDCE_1 (Q, C, CE, CLR, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input CLR ;
input D ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDCE_1 ####

//#### BEGIN MODULE DEFINITION FOR :FDCP ###
module FDCP (Q, C, CLR, D, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CLR ;
input D ;
input PRE ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDCP ####

//#### BEGIN MODULE DEFINITION FOR :FDCPE ###
module FDCPE (Q, C, CE, CLR, D, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input CLR ;
input D ;
input PRE ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDCPE ####

//#### BEGIN MODULE DEFINITION FOR :FDCPE_1 ###
module FDCPE_1 (Q, C, CE, CLR, D, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input CLR ;
input D ;
input PRE ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDCPE_1 ####

//#### BEGIN MODULE DEFINITION FOR :FDCP_1 ###
module FDCP_1 (Q, C, CLR, D, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CLR ;
input D ;
input PRE ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDCP_1 ####

//#### BEGIN MODULE DEFINITION FOR :FDC_1 ###
module FDC_1 (Q, C, CLR, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CLR ;
input D ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDC_1 ####

//#### BEGIN MODULE DEFINITION FOR :FDDRCPE ###
module FDDRCPE (Q, C0, C1, CE, CLR, D0, D1, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C0 ;
input C1 ;
input CE ;
input CLR ;
input D0 ;
input D1 ;
input PRE ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDDRCPE ####

//#### BEGIN MODULE DEFINITION FOR :FDDRRSE ###
module FDDRRSE (Q, C0, C1, CE, D0, D1, R, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C0 ;
input C1 ;
input CE ;
input D0 ;
input D1 ;
input R ;
input S ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDDRRSE ####

//#### BEGIN MODULE DEFINITION FOR :FDE ###
module FDE (Q, C, CE, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input D ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDE ####

//#### BEGIN MODULE DEFINITION FOR :FDE_1 ###
module FDE_1 (Q, C, CE, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input D ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDE_1 ####

//#### BEGIN MODULE DEFINITION FOR :FDP ###
module FDP (Q, C, D, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input D ;
input PRE ;
output Q ;
parameter INIT = 1'b1;
endmodule
//#### END MODULE DEFINITION FOR: FDP ####

//#### BEGIN MODULE DEFINITION FOR :FDPE ###
module FDPE (Q, C, CE, D, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input D ;
input PRE ;
output Q ;
parameter INIT = 1'b1;
endmodule
//#### END MODULE DEFINITION FOR: FDPE ####

//#### BEGIN MODULE DEFINITION FOR :FDPE_1 ###
module FDPE_1 (Q, C, CE, D, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input D ;
input PRE ;
output Q ;
parameter INIT = 1'b1;
endmodule
//#### END MODULE DEFINITION FOR: FDPE_1 ####

//#### BEGIN MODULE DEFINITION FOR :FDP_1 ###
module FDP_1 (Q, C, D, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input D ;
input PRE ;
output Q ;
parameter INIT = 1'b1;
endmodule
//#### END MODULE DEFINITION FOR: FDP_1 ####

//#### BEGIN MODULE DEFINITION FOR :FDR ###
module FDR (Q, C, D, R) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input D ;
input R ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDR ####

//#### BEGIN MODULE DEFINITION FOR :FDRE ###
module FDRE (Q, C, CE, D, R) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input D ;
input R ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDRE ####

//#### BEGIN MODULE DEFINITION FOR :FDRE_1 ###
module FDRE_1 (Q, C, CE, D, R) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input D ;
input R ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDRE_1 ####

//#### BEGIN MODULE DEFINITION FOR :FDRS ###
module FDRS (Q, C, D, R, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input D ;
input R ;
input S ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDRS ####

//#### BEGIN MODULE DEFINITION FOR :FDRSE ###
module FDRSE (Q, C, CE, D, R, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input D ;
input R ;
input S ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDRSE ####

//#### BEGIN MODULE DEFINITION FOR :FDRSE_1 ###
module FDRSE_1 (Q, C, CE, D, R, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input D ;
input R ;
input S ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDRSE_1 ####

//#### BEGIN MODULE DEFINITION FOR :FDRS_1 ###
module FDRS_1 (Q, C, D, R, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input D ;
input R ;
input S ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDRS_1 ####

//#### BEGIN MODULE DEFINITION FOR :FDR_1 ###
module FDR_1 (Q, C, D, R) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input D ;
input R ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FDR_1 ####

//#### BEGIN MODULE DEFINITION FOR :FDS ###
module FDS (Q, C, D, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input D ;
input S ;
output Q ;
parameter INIT = 1'b1;
endmodule
//#### END MODULE DEFINITION FOR: FDS ####

//#### BEGIN MODULE DEFINITION FOR :FDSE ###
module FDSE (Q, C, CE, D, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input D ;
input S ;
output Q ;
parameter INIT = 1'b1;
endmodule
//#### END MODULE DEFINITION FOR: FDSE ####

//#### BEGIN MODULE DEFINITION FOR :FDSE_1 ###
module FDSE_1 (Q, C, CE, D, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input D ;
input S ;
output Q ;
parameter INIT = 1'b1;
endmodule
//#### END MODULE DEFINITION FOR: FDSE_1 ####

//#### BEGIN MODULE DEFINITION FOR :FDS_1 ###
module FDS_1 (Q, C, D, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input D ;
input S ;
output Q ;
parameter INIT = 1'b1;
endmodule
//#### END MODULE DEFINITION FOR: FDS_1 ####

//#### BEGIN MODULE DEFINITION FOR :FD_1 ###
module FD_1 (Q, C, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input D ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: FD_1 ####

//#### BEGIN MODULE DEFINITION FOR :FIFO16 ###
module FIFO16 (ALMOSTEMPTY, ALMOSTFULL, DO, DOP, EMPTY, FULL, RDCOUNT, RDERR, WRCOUNT, WRERR, DI, DIP, RDCLK, RDEN, RST, WRCLK, WREN
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [31:0] DI ;
input [3:0] DIP ;
input RDCLK ;
input RDEN ;
input RST ;
input WRCLK ;
input WREN ;
output ALMOSTEMPTY ;
output ALMOSTFULL ;
output [31:0] DO ;
output [3:0] DOP ;
output EMPTY ;
output FULL ;
output [11:0] RDCOUNT ;
output RDERR ;
output [11:0] WRCOUNT ;
output WRERR ;
parameter ALMOST_FULL_OFFSET = 12'h080;
parameter ALMOST_EMPTY_OFFSET = 12'h080;
parameter DATA_WIDTH = 36;
parameter FIRST_WORD_FALL_THROUGH = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: FIFO16 ####

//#### BEGIN MODULE DEFINITION FOR :FIFO18 ###
module FIFO18 (ALMOSTEMPTY, ALMOSTFULL, DO, DOP, EMPTY, FULL, RDCOUNT, RDERR, WRCOUNT, WRERR,
	       DI, DIP, RDCLK, RDEN, RST, WRCLK, WREN) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [15:0] DI ;
input [1:0] DIP ;
input RDCLK ;
input RDEN ;
input RST ;
input WRCLK ;
input WREN ;
output ALMOSTEMPTY ;
output ALMOSTFULL ;
output [15:0] DO ;
output [1:0] DOP ;
output EMPTY ;
output FULL ;
output [11:0] RDCOUNT ;
output RDERR ;
output [11:0] WRCOUNT ;
output WRERR ;
parameter ALMOST_EMPTY_OFFSET = 12'h080;
parameter ALMOST_FULL_OFFSET = 12'h080;
parameter DATA_WIDTH = 4;
parameter DO_REG = 1;
parameter EN_SYN = "FALSE";
parameter FIRST_WORD_FALL_THROUGH = "FALSE";
parameter SIM_MODE = "SAFE";
endmodule
//#### END MODULE DEFINITION FOR: FIFO18 ####

//#### BEGIN MODULE DEFINITION FOR :FIFO18E1 ###
module FIFO18E1 (ALMOSTEMPTY, ALMOSTFULL, DO, DOP, EMPTY, FULL, RDCOUNT, RDERR, WRCOUNT, WRERR,
	       DI, DIP, RDCLK, RDEN, REGCE, RST, RSTREG, WRCLK, WREN) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [31:0] DI ;
input [3:0] DIP ;
input RDCLK ;
input RDEN ;
input REGCE ;
input RST ;
input RSTREG ;
input WRCLK ;
input WREN ;
output ALMOSTEMPTY ;
output ALMOSTFULL ;
output [31:0] DO ;
output [3:0] DOP ;
output EMPTY ;
output FULL ;
output [11:0] RDCOUNT ;
output RDERR ;
output [11:0] WRCOUNT ;
output WRERR ;
parameter ALMOST_EMPTY_OFFSET = 13'h0080;
parameter ALMOST_FULL_OFFSET = 13'h0080;
parameter DATA_WIDTH = 4;
parameter DO_REG = 1;
parameter EN_SYN = "FALSE";
parameter FIFO_MODE = "FIFO18";
parameter FIRST_WORD_FALL_THROUGH = "FALSE";
parameter INIT = 36'h0;
parameter SIM_DEVICE = "VIRTEX6";
parameter SRVAL = 36'h0;
endmodule
//#### END MODULE DEFINITION FOR: FIFO18E1 ####

//#### BEGIN MODULE DEFINITION FOR :FIFO18_36 ###
module FIFO18_36 (ALMOSTEMPTY, ALMOSTFULL, DO, DOP, EMPTY, FULL, RDCOUNT, RDERR, WRCOUNT, WRERR,
		  DI, DIP, RDCLK, RDEN, RST, WRCLK, WREN) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [31:0] DI ;
input [3:0] DIP ;
input RDCLK ;
input RDEN ;
input RST ;
input WRCLK ;
input WREN ;
output ALMOSTEMPTY ;
output ALMOSTFULL ;
output [31:0] DO ;
output [3:0] DOP ;
output EMPTY ;
output FULL ;
output [8:0] RDCOUNT ;
output RDERR ;
output [8:0] WRCOUNT ;
output WRERR ;
parameter ALMOST_EMPTY_OFFSET = 9'h080;
parameter ALMOST_FULL_OFFSET = 9'h080;
parameter DO_REG = 1;
parameter EN_SYN = "FALSE";
parameter FIRST_WORD_FALL_THROUGH = "FALSE";
parameter SIM_MODE = "SAFE";
endmodule
//#### END MODULE DEFINITION FOR: FIFO18_36 ####

//#### BEGIN MODULE DEFINITION FOR :FIFO36 ###
module FIFO36 (ALMOSTEMPTY, ALMOSTFULL, DO, DOP, EMPTY, FULL, RDCOUNT, RDERR, WRCOUNT, WRERR,
	       DI, DIP, RDCLK, RDEN, RST, WRCLK, WREN) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [31:0] DI ;
input [3:0] DIP ;
input RDCLK ;
input RDEN ;
input RST ;
input WRCLK ;
input WREN ;
output ALMOSTEMPTY ;
output ALMOSTFULL ;
output [31:0] DO ;
output [3:0] DOP ;
output EMPTY ;
output FULL ;
output [12:0] RDCOUNT ;
output RDERR ;
output [12:0] WRCOUNT ;
output WRERR ;
parameter ALMOST_EMPTY_OFFSET = 13'h0080;
parameter ALMOST_FULL_OFFSET = 13'h0080;
parameter DATA_WIDTH = 4;
parameter DO_REG = 1;
parameter EN_SYN = "FALSE";
parameter FIRST_WORD_FALL_THROUGH = "FALSE";
parameter SIM_MODE = "SAFE";
endmodule
//#### END MODULE DEFINITION FOR: FIFO36 ####

//#### BEGIN MODULE DEFINITION FOR :FIFO36E1 ###
module FIFO36E1 (ALMOSTEMPTY, ALMOSTFULL, DBITERR, DO, DOP, ECCPARITY, EMPTY, FULL, RDCOUNT, RDERR, SBITERR, WRCOUNT, WRERR,
	       DI, DIP, INJECTDBITERR, INJECTSBITERR, RDCLK, RDEN, REGCE, RST, RSTREG, WRCLK, WREN) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [63:0] DI ;
input [7:0] DIP ;
input INJECTDBITERR ;
input INJECTSBITERR ;
input RDCLK ;
input RDEN ;
input REGCE ;
input RST ;
input RSTREG ;
input WRCLK ;
input WREN ;
output ALMOSTEMPTY ;
output ALMOSTFULL ;
output DBITERR ;
output [63:0] DO ;
output [7:0] DOP ;
output [7:0] ECCPARITY ;
output EMPTY ;
output FULL ;
output [12:0] RDCOUNT ;
output RDERR ;
output SBITERR ;
output [12:0] WRCOUNT ;
output WRERR ;
parameter ALMOST_EMPTY_OFFSET = 13'h0080;
parameter ALMOST_FULL_OFFSET = 13'h0080;
parameter DATA_WIDTH = 4;
parameter DO_REG = 1;
parameter EN_ECC_READ = "FALSE";
parameter EN_ECC_WRITE = "FALSE";
parameter EN_SYN = "FALSE";
parameter FIFO_MODE = "FIFO36";
parameter FIRST_WORD_FALL_THROUGH = "FALSE";
parameter INIT = 72'h0;
parameter SIM_DEVICE = "VIRTEX6";
parameter SRVAL = 72'h0;
endmodule
//#### END MODULE DEFINITION FOR: FIFO36E1 ####

//#### BEGIN MODULE DEFINITION FOR :FIFO36_72 ###
module FIFO36_72 (ALMOSTEMPTY, ALMOSTFULL, DBITERR, DO, DOP, ECCPARITY, EMPTY, FULL, RDCOUNT, RDERR, SBITERR, WRCOUNT, WRERR,
	       DI, DIP, RDCLK, RDEN, RST, WRCLK, WREN) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [63:0] DI ;
input [7:0] DIP ;
input RDCLK ;
input RDEN ;
input RST ;
input WRCLK ;
input WREN ;
output ALMOSTEMPTY ;
output ALMOSTFULL ;
output DBITERR ;
output [63:0] DO ;
output [7:0] DOP ;
output [7:0] ECCPARITY ;
output EMPTY ;
output FULL ;
output [8:0] RDCOUNT ;
output RDERR ;
output SBITERR ;
output [8:0] WRCOUNT ;
output WRERR ;
parameter ALMOST_EMPTY_OFFSET = 9'h080;
parameter ALMOST_FULL_OFFSET = 9'h080;
parameter DO_REG = 1;
parameter EN_ECC_WRITE = "FALSE";
parameter EN_ECC_READ = "FALSE";
parameter EN_SYN = "FALSE";
parameter FIRST_WORD_FALL_THROUGH = "FALSE";
parameter SIM_MODE = "SAFE";
endmodule
//#### END MODULE DEFINITION FOR: FIFO36_72 ####

//#### BEGIN MODULE DEFINITION FOR :FIFO36_72_EXP ###
module FIFO36_72_EXP (ALMOSTEMPTY, ALMOSTFULL, DBITERR, DO, DOP, ECCPARITY, EMPTY, FULL, RDCOUNT, RDERR, SBITERR, WRCOUNT, WRERR,
		      DI, DIP, RDCLKL, RDCLKU, RDEN, RDRCLKL, RDRCLKU, RST, WRCLKL, WRCLKU, WREN) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [63:0] DI ;
input [7:0] DIP ;
input RDCLKL ;
input RDCLKU ;
input RDEN ;
input RDRCLKL ;
input RDRCLKU ;
input RST ;
input WRCLKL ;
input WRCLKU ;
input WREN ;
output ALMOSTEMPTY ;
output ALMOSTFULL ;
output DBITERR ;
output [63:0] DO ;
output [7:0] DOP ;
output [7:0] ECCPARITY ;
output EMPTY ;
output FULL ;
output [12:0] RDCOUNT ;
output RDERR ;
output SBITERR ;
output [12:0] WRCOUNT ;
output WRERR ;
parameter ALMOST_EMPTY_OFFSET = 9'h080;
parameter ALMOST_FULL_OFFSET = 9'h080;
parameter DO_REG = 1;
parameter EN_ECC_WRITE = "FALSE";
parameter EN_ECC_READ = "FALSE";
parameter EN_SYN = "FALSE";
parameter FIRST_WORD_FALL_THROUGH = "FALSE";
parameter SIM_MODE = "SAFE";
endmodule
//#### END MODULE DEFINITION FOR: FIFO36_72_EXP ####

//#### BEGIN MODULE DEFINITION FOR :FIFO36_EXP ###
module FIFO36_EXP (ALMOSTEMPTY, ALMOSTFULL, DO, DOP, EMPTY, FULL, RDCOUNT, RDERR, WRCOUNT, WRERR,
	       DI, DIP, RDCLKL, RDCLKU, RDEN, RDRCLKL, RDRCLKU, RST, WRCLKL, WRCLKU, WREN) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [31:0] DI ;
input [3:0] DIP ;
input RDCLKL ;
input RDCLKU ;
input RDEN ;
input RDRCLKL ;
input RDRCLKU ;
input RST ;
input WRCLKL ;
input WRCLKU ;
input WREN ;
output ALMOSTEMPTY ;
output ALMOSTFULL ;
output [31:0] DO ;
output [3:0] DOP ;
output EMPTY ;
output FULL ;
output [12:0] RDCOUNT ;
output RDERR ;
output [12:0] WRCOUNT ;
output WRERR ;
parameter ALMOST_EMPTY_OFFSET = 13'h0080;
parameter ALMOST_FULL_OFFSET = 13'h0080;
parameter DATA_WIDTH = 4;
parameter DO_REG = 1;
parameter EN_SYN = "FALSE";
parameter FIRST_WORD_FALL_THROUGH = "FALSE";
parameter SIM_MODE = "SAFE";
endmodule
//#### END MODULE DEFINITION FOR: FIFO36_EXP ####

//#### BEGIN MODULE DEFINITION FOR :FMAP ###
module FMAP (I1, I2, I3, I4, O) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
input O ;
endmodule
//#### END MODULE DEFINITION FOR: FMAP ####

//#### BEGIN MODULE DEFINITION FOR :FRAME_ECCE2 ###
module FRAME_ECCE2 (
  CRCERROR,
  ECCERROR,
  ECCERRORSINGLE,
  FAR,
  SYNBIT,
  SYNDROME,
  SYNDROMEVALID,
  SYNWORD
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
output CRCERROR ;
output ECCERROR ;
output ECCERRORSINGLE ;
output SYNDROMEVALID ;
output [12:0] SYNDROME ;
output [25:0] FAR ;
output [4:0] SYNBIT ;
output [6:0] SYNWORD ;
parameter FARSRC = "EFAR";
parameter FRAME_RBT_IN_FILENAME = "NONE";
endmodule
//#### END MODULE DEFINITION FOR: FRAME_ECCE2 ####

//#### BEGIN MODULE DEFINITION FOR :FRAME_ECC_VIRTEX4 ###
module FRAME_ECC_VIRTEX4 (ERROR, SYNDROME, SYNDROMEVALID) /* synthesis syn_black_box  syn_lib_cell=1
 */;
output ERROR ;
output [11:0] SYNDROME ;
output SYNDROMEVALID ;
endmodule
//#### END MODULE DEFINITION FOR: FRAME_ECC_VIRTEX4 ####

//#### BEGIN MODULE DEFINITION FOR :FRAME_ECC_VIRTEX5 ###
module FRAME_ECC_VIRTEX5 (
	CRCERROR,
	ECCERROR,
	SYNDROME,
	SYNDROMEVALID
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
output CRCERROR ;
output ECCERROR ;
output SYNDROMEVALID ;
output [11:0] SYNDROME ;
endmodule
//#### END MODULE DEFINITION FOR: FRAME_ECC_VIRTEX5 ####

//#### BEGIN MODULE DEFINITION FOR :FRAME_ECC_VIRTEX6 ###
module FRAME_ECC_VIRTEX6 (
  CRCERROR,
  ECCERROR,
  ECCERRORSINGLE,
  FAR,
  SYNBIT,
  SYNDROME,
  SYNDROMEVALID,
  SYNWORD
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
output CRCERROR ;
output ECCERROR ;
output ECCERRORSINGLE ;
output SYNDROMEVALID ;
output [12:0] SYNDROME ;
output [23:0] FAR ;
output [4:0] SYNBIT ;
output [6:0] SYNWORD ;
parameter FARSRC = "EFAR";
parameter FRAME_RBT_IN_FILENAME = "NONE";
endmodule
//#### END MODULE DEFINITION FOR: FRAME_ECC_VIRTEX6 ####

//#### BEGIN MODULE DEFINITION FOR :GND ###
module GND(G) /* synthesis syn_black_box  syn_lib_cell=1
 .noprune=1
 */;
output G ;
endmodule
//#### END MODULE DEFINITION FOR: GND ####

//#### BEGIN MODULE DEFINITION FOR :GT11 ###
module GT11 (
	CHBONDO,
	COMBUSOUT,
	DO,
	DRDY,
	RXBUFERR,
	RXCALFAIL,
	RXCHARISCOMMA,
	RXCHARISK,
	RXCOMMADET,
	RXCRCOUT,
	RXCYCLELIMIT,
	RXDATA,
	RXDISPERR,
	RXLOCK,
	RXLOSSOFSYNC,
	RXMCLK,
	RXNOTINTABLE,
	RXPCSHCLKOUT,
	RXREALIGN,
	RXRECCLK1,
	RXRECCLK2,
	RXRUNDISP,
	RXSIGDET,
	RXSTATUS,
	TX1N,
	TX1P,
	TXBUFERR,
	TXCALFAIL,
	TXCRCOUT,
	TXCYCLELIMIT,
	TXKERR,
	TXLOCK,
	TXOUTCLK1,
	TXOUTCLK2,
	TXPCSHCLKOUT,
	TXRUNDISP,
	CHBONDI,
	COMBUSIN,
	DADDR,
	DCLK,
	DEN,
	DI,
	DWE,
	ENCHANSYNC,
	ENMCOMMAALIGN,
	ENPCOMMAALIGN,
	GREFCLK,
	LOOPBACK,
	POWERDOWN,
	REFCLK1,
	REFCLK2,
	RX1N,
	RX1P,
	RXBLOCKSYNC64B66BUSE,
	RXCLKSTABLE,
	RXCOMMADETUSE,
	RXCRCCLK,
	RXCRCDATAVALID,
	RXCRCDATAWIDTH,
	RXCRCIN,
	RXCRCINIT,
	RXCRCINTCLK,
	RXCRCPD,
	RXCRCRESET,
	RXDATAWIDTH,
	RXDEC64B66BUSE,
	RXDEC8B10BUSE,
	RXDESCRAM64B66BUSE,
	RXIGNOREBTF,
	RXINTDATAWIDTH,
	RXPMARESET,
	RXPOLARITY,
	RXRESET,
	RXSLIDE,
	RXSYNC,
	RXUSRCLK,
	RXUSRCLK2,
	TXBYPASS8B10B,
	TXCHARDISPMODE,
	TXCHARDISPVAL,
	TXCHARISK,
	TXCLKSTABLE,
	TXCRCCLK,
	TXCRCDATAVALID,
	TXCRCDATAWIDTH,
	TXCRCIN,
	TXCRCINIT,
	TXCRCINTCLK,
	TXCRCPD,
	TXCRCRESET,
	TXDATA,
	TXDATAWIDTH,
	TXENC64B66BUSE,
	TXENC8B10BUSE,
	TXENOOB,
	TXGEARBOX64B66BUSE,
	TXINHIBIT,
	TXINTDATAWIDTH,
	TXPMARESET,
	TXPOLARITY,
	TXRESET,
	TXSCRAM64B66BUSE,
	TXSYNC,
	TXUSRCLK,
	TXUSRCLK2
) /* synthesis syn_black_box  syn_lib_cell=1
 black_box_pad_pin="RX1N,RX1P,TX1N,TX1P"
 */;
input DCLK ;
input DEN ;
input DWE ;
input ENCHANSYNC ;
input ENMCOMMAALIGN ;
input ENPCOMMAALIGN ;
input GREFCLK ;
input POWERDOWN ;
input REFCLK1 ;
input REFCLK2 ;
input RX1N ;
input RX1P ;
input RXBLOCKSYNC64B66BUSE ;
input RXCLKSTABLE ;
input RXCOMMADETUSE ;
input RXCRCCLK ;
input RXCRCDATAVALID ;
input RXCRCINIT ;
input RXCRCINTCLK ;
input RXCRCPD ;
input RXCRCRESET ;
input RXDEC64B66BUSE ;
input RXDEC8B10BUSE ;
input RXDESCRAM64B66BUSE ;
input RXIGNOREBTF ;
input RXPMARESET ;
input RXPOLARITY ;
input RXRESET ;
input RXSLIDE ;
input RXSYNC ;
input RXUSRCLK2 ;
input RXUSRCLK ;
input TXCLKSTABLE ;
input TXCRCCLK ;
input TXCRCDATAVALID ;
input TXCRCINIT ;
input TXCRCINTCLK ;
input TXCRCPD ;
input TXCRCRESET ;
input TXENC64B66BUSE ;
input TXENC8B10BUSE ;
input TXENOOB ;
input TXGEARBOX64B66BUSE ;
input TXINHIBIT ;
input TXPMARESET ;
input TXPOLARITY ;
input TXRESET ;
input TXSCRAM64B66BUSE ;
input TXSYNC ;
input TXUSRCLK2 ;
input TXUSRCLK ;
input [15:0] COMBUSIN ;
input [15:0] DI ;
input [1:0] LOOPBACK ;
input [1:0] RXDATAWIDTH ;
input [1:0] RXINTDATAWIDTH ;
input [1:0] TXDATAWIDTH ;
input [1:0] TXINTDATAWIDTH ;
input [2:0] RXCRCDATAWIDTH ;
input [2:0] TXCRCDATAWIDTH ;
input [4:0] CHBONDI ;
input [63:0] RXCRCIN ;
input [63:0] TXCRCIN ;
input [63:0] TXDATA ;
input [7:0] DADDR ;
input [7:0] TXBYPASS8B10B ;
input [7:0] TXCHARDISPMODE ;
input [7:0] TXCHARDISPVAL ;
input [7:0] TXCHARISK ;
output DRDY ;
output RXBUFERR ;
output RXCALFAIL ;
output RXCOMMADET ;
output RXCYCLELIMIT ;
output RXLOCK ;
output RXMCLK ;
output RXPCSHCLKOUT ;
output RXREALIGN ;
output RXRECCLK1 ;
output RXRECCLK2 ;
output RXSIGDET ;
output TX1N ;
output TX1P ;
output TXBUFERR ;
output TXCALFAIL ;
output TXCYCLELIMIT ;
output TXLOCK ;
output TXOUTCLK1 ;
output TXOUTCLK2 ;
output TXPCSHCLKOUT ;
output [15:0] COMBUSOUT ;
output [15:0] DO ;
output [1:0] RXLOSSOFSYNC ;
output [31:0] RXCRCOUT ;
output [31:0] TXCRCOUT ;
output [4:0] CHBONDO ;
output [5:0] RXSTATUS ;
output [63:0] RXDATA ;
output [7:0] RXCHARISCOMMA ;
output [7:0] RXCHARISK ;
output [7:0] RXDISPERR ;
output [7:0] RXNOTINTABLE ;
output [7:0] RXRUNDISP ;
output [7:0] TXKERR ;
output [7:0] TXRUNDISP ;
parameter BANDGAPSEL = "FALSE";
parameter BIASRESSEL = "FALSE";
parameter CCCB_ARBITRATOR_DISABLE = "FALSE";
parameter CHAN_BOND_MODE = "NONE";
parameter CHAN_BOND_ONE_SHOT = "FALSE";
parameter CHAN_BOND_SEQ_1_1 = 11'b00000000000;
parameter CHAN_BOND_SEQ_1_2 = 11'b00000000000;
parameter CHAN_BOND_SEQ_1_3 = 11'b00000000000;
parameter CHAN_BOND_SEQ_1_4 = 11'b00000000000;
parameter CHAN_BOND_SEQ_1_MASK = 4'b1110;
parameter CHAN_BOND_SEQ_2_1 = 11'b00000000000;
parameter CHAN_BOND_SEQ_2_2 = 11'b00000000000;
parameter CHAN_BOND_SEQ_2_3 = 11'b00000000000;
parameter CHAN_BOND_SEQ_2_4 = 11'b00000000000;
parameter CHAN_BOND_SEQ_2_MASK = 4'b1110;
parameter CHAN_BOND_SEQ_2_USE = "FALSE";
parameter CLK_CORRECT_USE = "FALSE";
parameter CLK_COR_8B10B_DE = "FALSE";
parameter CLK_COR_SEQ_1_1 = 11'b00000000000;
parameter CLK_COR_SEQ_1_2 = 11'b00000000000;
parameter CLK_COR_SEQ_1_3 = 11'b00000000000;
parameter CLK_COR_SEQ_1_4 = 11'b00000000000;
parameter CLK_COR_SEQ_1_MASK = 4'b1110;
parameter CLK_COR_SEQ_2_1 = 11'b00000000000;
parameter CLK_COR_SEQ_2_2 = 11'b00000000000;
parameter CLK_COR_SEQ_2_3 = 11'b00000000000;
parameter CLK_COR_SEQ_2_4 = 11'b00000000000;
parameter CLK_COR_SEQ_2_MASK = 4'b1110;
parameter CLK_COR_SEQ_2_USE = "FALSE";
parameter CLK_COR_SEQ_DROP = "FALSE";
parameter COMMA32 = "FALSE";
parameter COMMA_10B_MASK = 10'h3FF;
parameter CYCLE_LIMIT_SEL = 2'b00;
parameter DCDR_FILTER = 3'b010;
parameter DEC_MCOMMA_DETECT = "TRUE";
parameter DEC_PCOMMA_DETECT = "TRUE";
parameter DEC_VALID_COMMA_ONLY = "TRUE";
parameter DIGRX_FWDCLK = 2'b00;
parameter DIGRX_SYNC_MODE = "FALSE";
parameter ENABLE_DCDR = "FALSE";
parameter FDET_HYS_CAL = 3'b010;
parameter FDET_HYS_SEL = 3'b100;
parameter FDET_LCK_CAL = 3'b100;
parameter FDET_LCK_SEL = 3'b001;
parameter GT11_MODE = "DONT_CARE";
parameter IREFBIASMODE = 2'b11;
parameter LOOPCAL_WAIT = 2'b00;
parameter MCOMMA_32B_VALUE = 32'h00000000;
parameter MCOMMA_DETECT = "TRUE";
parameter OPPOSITE_SELECT = "FALSE";
parameter PCOMMA_32B_VALUE = 32'h00000000;
parameter PCOMMA_DETECT = "TRUE";
parameter PCS_BIT_SLIP = "FALSE";
parameter PMACLKENABLE = "TRUE";
parameter PMACOREPWRENABLE = "TRUE";
parameter PMAIREFTRIM = 4'b0111;
parameter PMAVBGCTRL = 5'b00000;
parameter PMAVREFTRIM = 4'b0111;
parameter PMA_BIT_SLIP = "FALSE";
parameter POWER_ENABLE = "TRUE";
parameter REPEATER = "FALSE";
parameter RXACTST = "FALSE";
parameter RXAFEEQ = 9'b000000000;
parameter RXAFEPD = "FALSE";
parameter RXAFETST = "FALSE";
parameter RXAPD = "FALSE";
parameter RXAREGCTRL = 5'b00000;
parameter RXASYNCDIVIDE = 2'b11;
parameter RXBY_32 = "FALSE";
parameter RXCDRLOS = 6'b000000;
parameter RXCLK0_FORCE_PMACLK = "FALSE";
parameter RXCLKMODE = 6'b110001;
parameter RXCLMODE = 2'b00;
parameter RXCMADJ = 2'b01;
parameter RXCPSEL = "TRUE";
parameter RXCPTST = "FALSE";
parameter RXCRCCLOCKDOUBLE = "FALSE";
parameter RXCRCENABLE = "FALSE";
parameter RXCRCINITVAL = 32'h00000000;
parameter RXCRCINVERTGEN = "FALSE";
parameter RXCRCSAMECLOCK = "FALSE";
parameter RXCTRL1 = 10'h200;
parameter RXCYCLE_LIMIT_SEL = 2'b00;
parameter RXDATA_SEL = 2'b00;
parameter RXDCCOUPLE = "FALSE";
parameter RXDIGRESET = "FALSE";
parameter RXDIGRX = "FALSE";
parameter RXEQ = 64'h4000000000000000;
parameter RXFDCAL_CLOCK_DIVIDE = "NONE";
parameter RXFDET_HYS_CAL = 3'b010;
parameter RXFDET_HYS_SEL = 3'b100;
parameter RXFDET_LCK_CAL = 3'b100;
parameter RXFDET_LCK_SEL = 3'b001;
parameter RXFECONTROL1 = 2'b00;
parameter RXFECONTROL2 = 3'b000;
parameter RXFETUNE = 2'b01;
parameter RXLB = "FALSE";
parameter RXLKADJ = 5'b00000;
parameter RXLKAPD = "FALSE";
parameter RXLOOPCAL_WAIT = 2'b00;
parameter RXLOOPFILT = 4'b0111;
parameter RXMODE = 6'b000000;
parameter RXPD = "FALSE";
parameter RXPDDTST = "TRUE";
parameter RXPMACLKSEL = "REFCLK1";
parameter RXRCPADJ = 3'b011;
parameter RXRCPPD = "FALSE";
parameter RXRECCLK1_USE_SYNC = "FALSE";
parameter RXRIBADJ = 2'b11;
parameter RXRPDPD = "FALSE";
parameter RXRSDPD = "FALSE";
parameter RXSLOWDOWN_CAL = 2'b00;
parameter RXTUNE = 13'h0000;
parameter RXVCODAC_INIT = 10'b1010000000;
parameter RXVCO_CTRL_ENABLE = "FALSE";
parameter RX_BUFFER_USE = "TRUE";
parameter RX_CLOCK_DIVIDER = 2'b00;
parameter SAMPLE_8X = "FALSE";
parameter SLOWDOWN_CAL = 2'b00;
parameter TXABPMACLKSEL = "REFCLK1";
parameter TXAPD = "FALSE";
parameter TXAREFBIASSEL = "TRUE";
parameter TXASYNCDIVIDE = 2'b11;
parameter TXCLK0_FORCE_PMACLK = "FALSE";
parameter TXCLKMODE = 4'b1001;
parameter TXCLMODE = 2'b00;
parameter TXCPSEL = "TRUE";
parameter TXCRCCLOCKDOUBLE = "FALSE";
parameter TXCRCENABLE = "FALSE";
parameter TXCRCINITVAL = 32'h00000000;
parameter TXCRCINVERTGEN = "FALSE";
parameter TXCRCSAMECLOCK = "FALSE";
parameter TXCTRL1 = 10'h200;
parameter TXDATA_SEL = 2'b00;
parameter TXDAT_PRDRV_DAC = 3'b111;
parameter TXDAT_TAP_DAC = 5'b10110;
parameter TXDIGPD = "FALSE";
parameter TXFDCAL_CLOCK_DIVIDE = "NONE";
parameter TXHIGHSIGNALEN = "TRUE";
parameter TXLOOPFILT = 4'b0111;
parameter TXLVLSHFTPD = "FALSE";
parameter TXOUTCLK1_USE_SYNC = "FALSE";
parameter TXPD = "FALSE";
parameter TXPHASESEL = "FALSE";
parameter TXPOST_PRDRV_DAC = 3'b111;
parameter TXPOST_TAP_DAC = 5'b01110;
parameter TXPOST_TAP_PD = "TRUE";
parameter TXPRE_PRDRV_DAC = 3'b111;
parameter TXPRE_TAP_DAC = 5'b00000;
parameter TXPRE_TAP_PD = "TRUE";
parameter TXSLEWRATE = "FALSE";
parameter TXTERMTRIM = 4'b1100;
parameter TXTUNE = 13'h0000;
parameter TX_BUFFER_USE = "TRUE";
parameter TX_CLOCK_DIVIDER = 2'b00;
parameter VCODAC_INIT = 10'b1010000000;
parameter VCO_CTRL_ENABLE = "FALSE";
parameter VREFBIASMODE = 2'b11;
parameter ALIGN_COMMA_WORD = 4;
parameter CHAN_BOND_LIMIT = 16;
parameter CHAN_BOND_SEQ_LEN = 1;
parameter CLK_COR_MAX_LAT = 48;
parameter CLK_COR_MIN_LAT = 36;
parameter CLK_COR_SEQ_LEN = 1;
parameter RXOUTDIV2SEL = 1;
parameter RXPLLNDIVSEL = 8;
parameter RXUSRDIVISOR = 1;
parameter SH_CNT_MAX = 64;
parameter SH_INVALID_CNT_MAX = 16;
parameter TXOUTDIV2SEL = 1;
parameter TXPLLNDIVSEL = 8;
endmodule
//#### END MODULE DEFINITION FOR: GT11 ####

//#### BEGIN MODULE DEFINITION FOR :GT11CLK ###
module GT11CLK (
	SYNCLK1OUT,
	SYNCLK2OUT,
	MGTCLKN,
	MGTCLKP,
	REFCLK,
	RXBCLK,
	SYNCLK1IN,
	SYNCLK2IN
) /* synthesis syn_black_box  syn_lib_cell=1
 black_box_pad_pin="MGTCLKN,MGTCLKP"
 */;
input MGTCLKN ;
input MGTCLKP ;
input REFCLK ;
input RXBCLK ;
input SYNCLK1IN ;
input SYNCLK2IN ;
output SYNCLK1OUT ;
output SYNCLK2OUT ;
parameter REFCLKSEL = "MGTCLK";
parameter SYNCLK1OUTEN = "ENABLE";
parameter SYNCLK2OUTEN = "DISABLE";
endmodule
//#### END MODULE DEFINITION FOR: GT11CLK ####

//#### BEGIN MODULE DEFINITION FOR :GT11CLK_MGT ###
module GT11CLK_MGT (
	SYNCLK1OUT,
	SYNCLK2OUT,
	MGTCLKN,
	MGTCLKP
) /* synthesis syn_black_box  syn_lib_cell=1
 black_box_pad_pin="MGTCLKN,MGTCLKP"
 */;
input MGTCLKN ;
input MGTCLKP ;
output SYNCLK1OUT ;
output SYNCLK2OUT ;
parameter SYNCLK1OUTEN = "ENABLE";
parameter SYNCLK2OUTEN = "DISABLE";
endmodule
//#### END MODULE DEFINITION FOR: GT11CLK_MGT ####

//#### BEGIN MODULE DEFINITION FOR :GT11_CUSTOM ###
module GT11_CUSTOM (
	CHBONDO,
	DO,
	DRDY,
	RXBUFERR,
	RXCALFAIL,
	RXCHARISCOMMA,
	RXCHARISK,
	RXCOMMADET,
	RXCRCOUT,
	RXCYCLELIMIT,
	RXDATA,
	RXDISPERR,
	RXLOCK,
	RXLOSSOFSYNC,
	RXMCLK,
	RXNOTINTABLE,
	RXPCSHCLKOUT,
	RXREALIGN,
	RXRECCLK1,
	RXRECCLK2,
	RXRUNDISP,
	RXSIGDET,
	RXSTATUS,
	TX1N,
	TX1P,
	TXBUFERR,
	TXCALFAIL,
	TXCRCOUT,
	TXCYCLELIMIT,
	TXKERR,
	TXLOCK,
	TXOUTCLK1,
	TXOUTCLK2,
	TXPCSHCLKOUT,
	TXRUNDISP,
	CHBONDI,
	DADDR,
	DCLK,
	DEN,
	DI,
	DWE,
	ENCHANSYNC,
	ENMCOMMAALIGN,
	ENPCOMMAALIGN,
	GREFCLK,
	LOOPBACK,
	POWERDOWN,
	REFCLK1,
	REFCLK2,
	RX1N,
	RX1P,
	RXBLOCKSYNC64B66BUSE,
	RXCLKSTABLE,
	RXCOMMADETUSE,
	RXCRCCLK,
	RXCRCDATAVALID,
	RXCRCDATAWIDTH,
	RXCRCIN,
	RXCRCINIT,
	RXCRCINTCLK,
	RXCRCPD,
	RXCRCRESET,
	RXDATAWIDTH,
	RXDEC64B66BUSE,
	RXDEC8B10BUSE,
	RXDESCRAM64B66BUSE,
	RXIGNOREBTF,
	RXINTDATAWIDTH,
	RXPMARESET,
	RXPOLARITY,
	RXRESET,
	RXSLIDE,
	RXSYNC,
	RXUSRCLK,
	RXUSRCLK2,
	TXBYPASS8B10B,
	TXCHARDISPMODE,
	TXCHARDISPVAL,
	TXCHARISK,
	TXCLKSTABLE,
	TXCRCCLK,
	TXCRCDATAVALID,
	TXCRCDATAWIDTH,
	TXCRCIN,
	TXCRCINIT,
	TXCRCINTCLK,
	TXCRCPD,
	TXCRCRESET,
	TXDATA,
	TXDATAWIDTH,
	TXENC64B66BUSE,
	TXENC8B10BUSE,
	TXENOOB,
	TXGEARBOX64B66BUSE,
	TXINHIBIT,
	TXINTDATAWIDTH,
	TXPMARESET,
	TXPOLARITY,
	TXRESET,
	TXSCRAM64B66BUSE,
	TXSYNC,
	TXUSRCLK,
	TXUSRCLK2
) /* synthesis syn_black_box  syn_lib_cell=1
 black_box_pad_pin="RX1N,RX1P,TX1N,TX1P"
 */;
input DCLK ;
input DEN ;
input DWE ;
input ENCHANSYNC ;
input ENMCOMMAALIGN ;
input ENPCOMMAALIGN ;
input GREFCLK ;
input POWERDOWN ;
input REFCLK1 ;
input REFCLK2 ;
input RX1N ;
input RX1P ;
input RXBLOCKSYNC64B66BUSE ;
input RXCLKSTABLE ;
input RXCOMMADETUSE ;
input RXCRCCLK ;
input RXCRCDATAVALID ;
input RXCRCINIT ;
input RXCRCINTCLK ;
input RXCRCPD ;
input RXCRCRESET ;
input RXDEC64B66BUSE ;
input RXDEC8B10BUSE ;
input RXDESCRAM64B66BUSE ;
input RXIGNOREBTF ;
input RXPMARESET ;
input RXPOLARITY ;
input RXRESET ;
input RXSLIDE ;
input RXSYNC ;
input RXUSRCLK2 ;
input RXUSRCLK ;
input TXCLKSTABLE ;
input TXCRCCLK ;
input TXCRCDATAVALID ;
input TXCRCINIT ;
input TXCRCINTCLK ;
input TXCRCPD ;
input TXCRCRESET ;
input TXENC64B66BUSE ;
input TXENC8B10BUSE ;
input TXENOOB ;
input TXGEARBOX64B66BUSE ;
input TXINHIBIT ;
input TXPMARESET ;
input TXPOLARITY ;
input TXRESET ;
input TXSCRAM64B66BUSE ;
input TXSYNC ;
input TXUSRCLK2 ;
input TXUSRCLK ;
input [15:0] DI ;
input [1:0] LOOPBACK ;
input [1:0] RXDATAWIDTH ;
input [1:0] RXINTDATAWIDTH ;
input [1:0] TXDATAWIDTH ;
input [1:0] TXINTDATAWIDTH ;
input [2:0] RXCRCDATAWIDTH ;
input [2:0] TXCRCDATAWIDTH ;
input [4:0] CHBONDI ;
input [63:0] RXCRCIN ;
input [63:0] TXCRCIN ;
input [63:0] TXDATA ;
input [7:0] DADDR ;
input [7:0] TXBYPASS8B10B ;
input [7:0] TXCHARDISPMODE ;
input [7:0] TXCHARDISPVAL ;
input [7:0] TXCHARISK ;
output DRDY ;
output RXBUFERR ;
output RXCALFAIL ;
output RXCOMMADET ;
output RXCYCLELIMIT ;
output RXLOCK ;
output RXMCLK ;
output RXPCSHCLKOUT ;
output RXREALIGN ;
output RXRECCLK1 ;
output RXRECCLK2 ;
output RXSIGDET ;
output TX1N ;
output TX1P ;
output TXBUFERR ;
output TXCALFAIL ;
output TXCYCLELIMIT ;
output TXLOCK ;
output TXOUTCLK1 ;
output TXOUTCLK2 ;
output TXPCSHCLKOUT ;
output [15:0] DO ;
output [1:0] RXLOSSOFSYNC ;
output [31:0] RXCRCOUT ;
output [31:0] TXCRCOUT ;
output [4:0] CHBONDO ;
output [5:0] RXSTATUS ;
output [63:0] RXDATA ;
output [7:0] RXCHARISCOMMA ;
output [7:0] RXCHARISK ;
output [7:0] RXDISPERR ;
output [7:0] RXNOTINTABLE ;
output [7:0] RXRUNDISP ;
output [7:0] TXKERR ;
output [7:0] TXRUNDISP ;
parameter BANDGAPSEL = "FALSE";
parameter BIASRESSEL = "FALSE";
parameter CCCB_ARBITRATOR_DISABLE = "FALSE";
parameter CHAN_BOND_MODE = "NONE";
parameter CHAN_BOND_ONE_SHOT = "FALSE";
parameter CHAN_BOND_SEQ_1_1 = 11'b00000000000;
parameter CHAN_BOND_SEQ_1_2 = 11'b00000000000;
parameter CHAN_BOND_SEQ_1_3 = 11'b00000000000;
parameter CHAN_BOND_SEQ_1_4 = 11'b00000000000;
parameter CHAN_BOND_SEQ_1_MASK = 4'b1110;
parameter CHAN_BOND_SEQ_2_1 = 11'b00000000000;
parameter CHAN_BOND_SEQ_2_2 = 11'b00000000000;
parameter CHAN_BOND_SEQ_2_3 = 11'b00000000000;
parameter CHAN_BOND_SEQ_2_4 = 11'b00000000000;
parameter CHAN_BOND_SEQ_2_MASK = 4'b1110;
parameter CHAN_BOND_SEQ_2_USE = "FALSE";
parameter CLK_CORRECT_USE = "FALSE";
parameter CLK_COR_8B10B_DE = "FALSE";
parameter CLK_COR_SEQ_1_1 = 11'b00000000000;
parameter CLK_COR_SEQ_1_2 = 11'b00000000000;
parameter CLK_COR_SEQ_1_3 = 11'b00000000000;
parameter CLK_COR_SEQ_1_4 = 11'b00000000000;
parameter CLK_COR_SEQ_1_MASK = 4'b1110;
parameter CLK_COR_SEQ_2_1 = 11'b00000000000;
parameter CLK_COR_SEQ_2_2 = 11'b00000000000;
parameter CLK_COR_SEQ_2_3 = 11'b00000000000;
parameter CLK_COR_SEQ_2_4 = 11'b00000000000;
parameter CLK_COR_SEQ_2_MASK = 4'b1110;
parameter CLK_COR_SEQ_2_USE = "FALSE";
parameter CLK_COR_SEQ_DROP = "FALSE";
parameter COMMA32 = "FALSE";
parameter COMMA_10B_MASK = 10'h3FF;
parameter CYCLE_LIMIT_SEL = 2'b00;
parameter DCDR_FILTER = 3'b010;
parameter DEC_MCOMMA_DETECT = "TRUE";
parameter DEC_PCOMMA_DETECT = "TRUE";
parameter DEC_VALID_COMMA_ONLY = "TRUE";
parameter DIGRX_FWDCLK = 2'b00;
parameter DIGRX_SYNC_MODE = "FALSE";
parameter ENABLE_DCDR = "FALSE";
parameter FDET_HYS_CAL = 3'b010;
parameter FDET_HYS_SEL = 3'b100;
parameter FDET_LCK_CAL = 3'b100;
parameter FDET_LCK_SEL = 3'b001;
parameter IREFBIASMODE = 2'b11;
parameter LOOPCAL_WAIT = 2'b00;
parameter MCOMMA_32B_VALUE = 32'h00000000;
parameter MCOMMA_DETECT = "TRUE";
parameter OPPOSITE_SELECT = "FALSE";
parameter PCOMMA_32B_VALUE = 32'h00000000;
parameter PCOMMA_DETECT = "TRUE";
parameter PCS_BIT_SLIP = "FALSE";
parameter PMACLKENABLE = "TRUE";
parameter PMACOREPWRENABLE = "TRUE";
parameter PMAIREFTRIM = 4'b0111;
parameter PMAVBGCTRL = 5'b00000;
parameter PMAVREFTRIM = 4'b0111;
parameter PMA_BIT_SLIP = "FALSE";
parameter POWER_ENABLE = "TRUE";
parameter REPEATER = "FALSE";
parameter RXACTST = "FALSE";
parameter RXAFEEQ = 9'b000000000;
parameter RXAFEPD = "FALSE";
parameter RXAFETST = "FALSE";
parameter RXAPD = "FALSE";
parameter RXAREGCTRL = 5'b00000;
parameter RXASYNCDIVIDE = 2'b11;
parameter RXBY_32 = "FALSE";
parameter RXCDRLOS = 6'b000000;
parameter RXCLK0_FORCE_PMACLK = "FALSE";
parameter RXCLKMODE = 6'b110001;
parameter RXCLMODE = 2'b00;
parameter RXCMADJ = 2'b01;
parameter RXCPSEL = "TRUE";
parameter RXCPTST = "FALSE";
parameter RXCRCCLOCKDOUBLE = "FALSE";
parameter RXCRCENABLE = "FALSE";
parameter RXCRCINITVAL = 32'h00000000;
parameter RXCRCINVERTGEN = "FALSE";
parameter RXCRCSAMECLOCK = "FALSE";
parameter RXCTRL1 = 10'h200;
parameter RXCYCLE_LIMIT_SEL = 2'b00;
parameter RXDATA_SEL = 2'b00;
parameter RXDCCOUPLE = "FALSE";
parameter RXDIGRESET = "FALSE";
parameter RXDIGRX = "FALSE";
parameter RXEQ = 64'h4000000000000000;
parameter RXFDCAL_CLOCK_DIVIDE = "NONE";
parameter RXFDET_HYS_CAL = 3'b010;
parameter RXFDET_HYS_SEL = 3'b100;
parameter RXFDET_LCK_CAL = 3'b100;
parameter RXFDET_LCK_SEL = 3'b001;
parameter RXFECONTROL1 = 2'b00;
parameter RXFECONTROL2 = 3'b000;
parameter RXFETUNE = 2'b01;
parameter RXLB = "FALSE";
parameter RXLKADJ = 5'b00000;
parameter RXLKAPD = "FALSE";
parameter RXLOOPCAL_WAIT = 2'b00;
parameter RXLOOPFILT = 4'b0111;
parameter RXMODE = 6'b000000;
parameter RXPD = "FALSE";
parameter RXPDDTST = "TRUE";
parameter RXPMACLKSEL = "REFCLK1";
parameter RXRCPADJ = 3'b011;
parameter RXRCPPD = "FALSE";
parameter RXRECCLK1_USE_SYNC = "FALSE";
parameter RXRIBADJ = 2'b11;
parameter RXRPDPD = "FALSE";
parameter RXRSDPD = "FALSE";
parameter RXSLOWDOWN_CAL = 2'b00;
parameter RXTUNE = 13'h0000;
parameter RXVCODAC_INIT = 10'b1010000000;
parameter RXVCO_CTRL_ENABLE = "FALSE";
parameter RX_BUFFER_USE = "TRUE";
parameter RX_CLOCK_DIVIDER = 2'b00;
parameter SAMPLE_8X = "FALSE";
parameter SLOWDOWN_CAL = 2'b00;
parameter TXABPMACLKSEL = "REFCLK1";
parameter TXAPD = "FALSE";
parameter TXAREFBIASSEL = "TRUE";
parameter TXASYNCDIVIDE = 2'b11;
parameter TXCLK0_FORCE_PMACLK = "FALSE";
parameter TXCLKMODE = 4'b1001;
parameter TXCLMODE = 2'b00;
parameter TXCPSEL = "TRUE";
parameter TXCRCCLOCKDOUBLE = "FALSE";
parameter TXCRCENABLE = "FALSE";
parameter TXCRCINITVAL = 32'h00000000;
parameter TXCRCINVERTGEN = "FALSE";
parameter TXCRCSAMECLOCK = "FALSE";
parameter TXCTRL1 = 10'h200;
parameter TXDATA_SEL = 2'b00;
parameter TXDAT_PRDRV_DAC = 3'b111;
parameter TXDAT_TAP_DAC = 5'b10110;
parameter TXDIGPD = "FALSE";
parameter TXFDCAL_CLOCK_DIVIDE = "NONE";
parameter TXHIGHSIGNALEN = "TRUE";
parameter TXLOOPFILT = 4'b0111;
parameter TXLVLSHFTPD = "FALSE";
parameter TXOUTCLK1_USE_SYNC = "FALSE";
parameter TXPD = "FALSE";
parameter TXPHASESEL = "FALSE";
parameter TXPOST_PRDRV_DAC = 3'b111;
parameter TXPOST_TAP_DAC = 5'b01110;
parameter TXPOST_TAP_PD = "TRUE";
parameter TXPRE_PRDRV_DAC = 3'b111;
parameter TXPRE_TAP_DAC = 5'b00000;
parameter TXPRE_TAP_PD = "TRUE";
parameter TXSLEWRATE = "FALSE";
parameter TXTERMTRIM = 4'b1100;
parameter TXTUNE = 13'h0000;
parameter TX_BUFFER_USE = "TRUE";
parameter TX_CLOCK_DIVIDER = 2'b00;
parameter VCODAC_INIT = 10'b1010000000;
parameter VCO_CTRL_ENABLE = "FALSE";
parameter VREFBIASMODE = 2'b11;
parameter ALIGN_COMMA_WORD = 4;
parameter CHAN_BOND_LIMIT = 16;
parameter CHAN_BOND_SEQ_LEN = 1;
parameter CLK_COR_MAX_LAT = 48;
parameter CLK_COR_MIN_LAT = 36;
parameter CLK_COR_SEQ_LEN = 1;
parameter RXOUTDIV2SEL = 1;
parameter RXPLLNDIVSEL = 8;
parameter RXUSRDIVISOR = 1;
parameter SH_CNT_MAX = 64;
parameter SH_INVALID_CNT_MAX = 16;
parameter TXOUTDIV2SEL = 1;
parameter TXPLLNDIVSEL = 8;
endmodule
//#### END MODULE DEFINITION FOR: GT11_CUSTOM ####

//#### BEGIN MODULE DEFINITION FOR :GT11_DUAL ###
module GT11_DUAL (
	CHBONDOA,
	CHBONDOB,
	DOA,
	DOB,
	DRDYA,
	DRDYB,
	RXBUFERRA,
	RXBUFERRB,
	RXCALFAILA,
	RXCALFAILB,
	RXCHARISCOMMAA,
	RXCHARISCOMMAB,
	RXCHARISKA,
	RXCHARISKB,
	RXCOMMADETA,
	RXCOMMADETB,
	RXCRCOUTA,
	RXCRCOUTB,
	RXCYCLELIMITA,
	RXCYCLELIMITB,
	RXDATAA,
	RXDATAB,
	RXDISPERRA,
	RXDISPERRB,
	RXLOCKA,
	RXLOCKB,
	RXLOSSOFSYNCA,
	RXLOSSOFSYNCB,
	RXMCLKA,
	RXMCLKB,
	RXNOTINTABLEA,
	RXNOTINTABLEB,
	RXPCSHCLKOUTA,
	RXPCSHCLKOUTB,
	RXREALIGNA,
	RXREALIGNB,
	RXRECCLK1A,
	RXRECCLK1B,
	RXRECCLK2A,
	RXRECCLK2B,
	RXRUNDISPA,
	RXRUNDISPB,
	RXSIGDETA,
	RXSIGDETB,
	RXSTATUSA,
	RXSTATUSB,
	TX1NA,
	TX1NB,
	TX1PA,
	TX1PB,
	TXBUFERRA,
	TXBUFERRB,
	TXCALFAILA,
	TXCALFAILB,
	TXCRCOUTA,
	TXCRCOUTB,
	TXCYCLELIMITA,
	TXCYCLELIMITB,
	TXKERRA,
	TXKERRB,
	TXLOCKA,
	TXLOCKB,
	TXOUTCLK1A,
	TXOUTCLK1B,
	TXOUTCLK2A,
	TXOUTCLK2B,
	TXPCSHCLKOUTA,
	TXPCSHCLKOUTB,
	TXRUNDISPA,
	TXRUNDISPB,
	CHBONDIA,
	CHBONDIB,
	DADDRA,
	DADDRB,
	DCLKA,
	DCLKB,
	DENA,
	DENB,
	DIA,
	DIB,
	DWEA,
	DWEB,
	ENCHANSYNCA,
	ENCHANSYNCB,
	ENMCOMMAALIGNA,
	ENMCOMMAALIGNB,
	ENPCOMMAALIGNA,
	ENPCOMMAALIGNB,
	GREFCLKA,
	GREFCLKB,
	LOOPBACKA,
	LOOPBACKB,
	POWERDOWNA,
	POWERDOWNB,
	REFCLK1A,
	REFCLK1B,
	REFCLK2A,
	REFCLK2B,
	RX1NA,
	RX1NB,
	RX1PA,
	RX1PB,
	RXBLOCKSYNC64B66BUSEA,
	RXBLOCKSYNC64B66BUSEB,
	RXCLKSTABLEA,
	RXCLKSTABLEB,
	RXCOMMADETUSEA,
	RXCOMMADETUSEB,
	RXCRCCLKA,
	RXCRCCLKB,
	RXCRCDATAVALIDA,
	RXCRCDATAVALIDB,
	RXCRCDATAWIDTHA,
	RXCRCDATAWIDTHB,
	RXCRCINA,
	RXCRCINB,
	RXCRCINITA,
	RXCRCINITB,
	RXCRCINTCLKA,
	RXCRCINTCLKB,
	RXCRCPDA,
	RXCRCPDB,
	RXCRCRESETA,
	RXCRCRESETB,
	RXDATAWIDTHA,
	RXDATAWIDTHB,
	RXDEC64B66BUSEA,
	RXDEC64B66BUSEB,
	RXDEC8B10BUSEA,
	RXDEC8B10BUSEB,
	RXDESCRAM64B66BUSEA,
	RXDESCRAM64B66BUSEB,
	RXIGNOREBTFA,
	RXIGNOREBTFB,
	RXINTDATAWIDTHA,
	RXINTDATAWIDTHB,
	RXPMARESETA,
	RXPMARESETB,
	RXPOLARITYA,
	RXPOLARITYB,
	RXRESETA,
	RXRESETB,
	RXSLIDEA,
	RXSLIDEB,
	RXSYNCA,
	RXSYNCB,
	RXUSRCLK2A,
	RXUSRCLK2B,
	RXUSRCLKA,
	RXUSRCLKB,
	TXBYPASS8B10BA,
	TXBYPASS8B10BB,
	TXCHARDISPMODEA,
	TXCHARDISPMODEB,
	TXCHARDISPVALA,
	TXCHARDISPVALB,
	TXCHARISKA,
	TXCHARISKB,
	TXCLKSTABLEA,
	TXCLKSTABLEB,
	TXCRCCLKA,
	TXCRCCLKB,
	TXCRCDATAVALIDA,
	TXCRCDATAVALIDB,
	TXCRCDATAWIDTHA,
	TXCRCDATAWIDTHB,
	TXCRCINA,
	TXCRCINB,
	TXCRCINITA,
	TXCRCINITB,
	TXCRCINTCLKA,
	TXCRCINTCLKB,
	TXCRCPDA,
	TXCRCPDB,
	TXCRCRESETA,
	TXCRCRESETB,
	TXDATAA,
	TXDATAB,
	TXDATAWIDTHA,
	TXDATAWIDTHB,
	TXENC64B66BUSEA,
	TXENC64B66BUSEB,
	TXENC8B10BUSEA,
	TXENC8B10BUSEB,
	TXENOOBA,
	TXENOOBB,
	TXGEARBOX64B66BUSEA,
	TXGEARBOX64B66BUSEB,
	TXINHIBITA,
	TXINHIBITB,
	TXINTDATAWIDTHA,
	TXINTDATAWIDTHB,
	TXPMARESETA,
	TXPMARESETB,
	TXPOLARITYA,
	TXPOLARITYB,
	TXRESETA,
	TXRESETB,
	TXSCRAM64B66BUSEA,
	TXSCRAM64B66BUSEB,
	TXSYNCA,
	TXSYNCB,
	TXUSRCLK2A,
	TXUSRCLK2B,
	TXUSRCLKA,
	TXUSRCLKB
) /* synthesis syn_black_box  syn_lib_cell=1
 black_box_pad_pin="RX1NA,RX1NB,RX1PA,RX1PB,TX1NA,TX1NB,TX1PA,TX1PB"
 */;
input DCLKA ;
input DCLKB ;
input DENA ;
input DENB ;
input DWEA ;
input DWEB ;
input ENCHANSYNCA ;
input ENCHANSYNCB ;
input ENMCOMMAALIGNA ;
input ENMCOMMAALIGNB ;
input ENPCOMMAALIGNA ;
input ENPCOMMAALIGNB ;
input GREFCLKA ;
input GREFCLKB ;
input POWERDOWNA ;
input POWERDOWNB ;
input REFCLK1A ;
input REFCLK1B ;
input REFCLK2A ;
input REFCLK2B ;
input RX1NA ;
input RX1NB ;
input RX1PA ;
input RX1PB ;
input RXBLOCKSYNC64B66BUSEA ;
input RXBLOCKSYNC64B66BUSEB ;
input RXCLKSTABLEA ;
input RXCLKSTABLEB ;
input RXCOMMADETUSEA ;
input RXCOMMADETUSEB ;
input RXCRCCLKA ;
input RXCRCCLKB ;
input RXCRCDATAVALIDA ;
input RXCRCDATAVALIDB ;
input RXCRCINITA ;
input RXCRCINITB ;
input RXCRCINTCLKA ;
input RXCRCINTCLKB ;
input RXCRCPDA ;
input RXCRCPDB ;
input RXCRCRESETA ;
input RXCRCRESETB ;
input RXDEC64B66BUSEA ;
input RXDEC64B66BUSEB ;
input RXDEC8B10BUSEA ;
input RXDEC8B10BUSEB ;
input RXDESCRAM64B66BUSEA ;
input RXDESCRAM64B66BUSEB ;
input RXIGNOREBTFA ;
input RXIGNOREBTFB ;
input RXPMARESETA ;
input RXPMARESETB ;
input RXPOLARITYA ;
input RXPOLARITYB ;
input RXRESETA ;
input RXRESETB ;
input RXSLIDEA ;
input RXSLIDEB ;
input RXSYNCA ;
input RXSYNCB ;
input RXUSRCLK2A ;
input RXUSRCLK2B ;
input RXUSRCLKA ;
input RXUSRCLKB ;
input TXCLKSTABLEA ;
input TXCLKSTABLEB ;
input TXCRCCLKA ;
input TXCRCCLKB ;
input TXCRCDATAVALIDA ;
input TXCRCDATAVALIDB ;
input TXCRCINITA ;
input TXCRCINITB ;
input TXCRCINTCLKA ;
input TXCRCINTCLKB ;
input TXCRCPDA ;
input TXCRCPDB ;
input TXCRCRESETA ;
input TXCRCRESETB ;
input TXENC64B66BUSEA ;
input TXENC64B66BUSEB ;
input TXENC8B10BUSEA ;
input TXENC8B10BUSEB ;
input TXENOOBA ;
input TXENOOBB ;
input TXGEARBOX64B66BUSEA ;
input TXGEARBOX64B66BUSEB ;
input TXINHIBITA ;
input TXINHIBITB ;
input TXPMARESETA ;
input TXPMARESETB ;
input TXPOLARITYA ;
input TXPOLARITYB ;
input TXRESETA ;
input TXRESETB ;
input TXSCRAM64B66BUSEA ;
input TXSCRAM64B66BUSEB ;
input TXSYNCA ;
input TXSYNCB ;
input TXUSRCLK2A ;
input TXUSRCLK2B ;
input TXUSRCLKA ;
input TXUSRCLKB ;
input [15:0] DIA ;
input [15:0] DIB ;
input [1:0] LOOPBACKA ;
input [1:0] LOOPBACKB ;
input [1:0] RXDATAWIDTHA ;
input [1:0] RXDATAWIDTHB ;
input [1:0] RXINTDATAWIDTHA ;
input [1:0] RXINTDATAWIDTHB ;
input [1:0] TXDATAWIDTHA ;
input [1:0] TXDATAWIDTHB ;
input [1:0] TXINTDATAWIDTHA ;
input [1:0] TXINTDATAWIDTHB ;
input [2:0] RXCRCDATAWIDTHA ;
input [2:0] RXCRCDATAWIDTHB ;
input [2:0] TXCRCDATAWIDTHA ;
input [2:0] TXCRCDATAWIDTHB ;
input [4:0] CHBONDIA ;
input [4:0] CHBONDIB ;
input [63:0] RXCRCINA ;
input [63:0] RXCRCINB ;
input [63:0] TXCRCINA ;
input [63:0] TXCRCINB ;
input [63:0] TXDATAA ;
input [63:0] TXDATAB ;
input [7:0] DADDRA ;
input [7:0] DADDRB ;
input [7:0] TXBYPASS8B10BA ;
input [7:0] TXBYPASS8B10BB ;
input [7:0] TXCHARDISPMODEA ;
input [7:0] TXCHARDISPMODEB ;
input [7:0] TXCHARDISPVALA ;
input [7:0] TXCHARDISPVALB ;
input [7:0] TXCHARISKA ;
input [7:0] TXCHARISKB ;
output DRDYA ;
output DRDYB ;
output RXBUFERRA ;
output RXBUFERRB ;
output RXCALFAILA ;
output RXCALFAILB ;
output RXCOMMADETA ;
output RXCOMMADETB ;
output RXCYCLELIMITA ;
output RXCYCLELIMITB ;
output RXLOCKA ;
output RXLOCKB ;
output RXMCLKA ;
output RXMCLKB ;
output RXPCSHCLKOUTA ;
output RXPCSHCLKOUTB ;
output RXREALIGNA ;
output RXREALIGNB ;
output RXRECCLK1A ;
output RXRECCLK1B ;
output RXRECCLK2A ;
output RXRECCLK2B ;
output RXSIGDETA ;
output RXSIGDETB ;
output TX1NA ;
output TX1NB ;
output TX1PA ;
output TX1PB ;
output TXBUFERRA ;
output TXBUFERRB ;
output TXCALFAILA ;
output TXCALFAILB ;
output TXCYCLELIMITA ;
output TXCYCLELIMITB ;
output TXLOCKA ;
output TXLOCKB ;
output TXOUTCLK1A ;
output TXOUTCLK1B ;
output TXOUTCLK2A ;
output TXOUTCLK2B ;
output TXPCSHCLKOUTA ;
output TXPCSHCLKOUTB ;
output [15:0] DOA ;
output [15:0] DOB ;
output [1:0] RXLOSSOFSYNCA ;
output [1:0] RXLOSSOFSYNCB ;
output [31:0] RXCRCOUTA ;
output [31:0] RXCRCOUTB ;
output [31:0] TXCRCOUTA ;
output [31:0] TXCRCOUTB ;
output [4:0] CHBONDOA ;
output [4:0] CHBONDOB ;
output [5:0] RXSTATUSA ;
output [5:0] RXSTATUSB ;
output [63:0] RXDATAA ;
output [63:0] RXDATAB ;
output [7:0] RXCHARISCOMMAA ;
output [7:0] RXCHARISCOMMAB ;
output [7:0] RXCHARISKA ;
output [7:0] RXCHARISKB ;
output [7:0] RXDISPERRA ;
output [7:0] RXDISPERRB ;
output [7:0] RXNOTINTABLEA ;
output [7:0] RXNOTINTABLEB ;
output [7:0] RXRUNDISPA ;
output [7:0] RXRUNDISPB ;
output [7:0] TXKERRA ;
output [7:0] TXKERRB ;
output [7:0] TXRUNDISPA ;
output [7:0] TXRUNDISPB ;
parameter BANDGAPSEL_A = "FALSE";
parameter BANDGAPSEL_B = "FALSE";
parameter BIASRESSEL_A = "FALSE";
parameter BIASRESSEL_B = "FALSE";
parameter CCCB_ARBITRATOR_DISABLE_A = "FALSE";
parameter CCCB_ARBITRATOR_DISABLE_B = "FALSE";
parameter CHAN_BOND_MODE_A = "NONE";
parameter CHAN_BOND_MODE_B = "NONE";
parameter CHAN_BOND_ONE_SHOT_A = "FALSE";
parameter CHAN_BOND_ONE_SHOT_B = "FALSE";
parameter CHAN_BOND_SEQ_1_1_A = 11'b00000000000;
parameter CHAN_BOND_SEQ_1_1_B = 11'b00000000000;
parameter CHAN_BOND_SEQ_1_2_A = 11'b00000000000;
parameter CHAN_BOND_SEQ_1_2_B = 11'b00000000000;
parameter CHAN_BOND_SEQ_1_3_A = 11'b00000000000;
parameter CHAN_BOND_SEQ_1_3_B = 11'b00000000000;
parameter CHAN_BOND_SEQ_1_4_A = 11'b00000000000;
parameter CHAN_BOND_SEQ_1_4_B = 11'b00000000000;
parameter CHAN_BOND_SEQ_1_MASK_A = 4'b1110;
parameter CHAN_BOND_SEQ_1_MASK_B = 4'b1110;
parameter CHAN_BOND_SEQ_2_1_A = 11'b00000000000;
parameter CHAN_BOND_SEQ_2_1_B = 11'b00000000000;
parameter CHAN_BOND_SEQ_2_2_A = 11'b00000000000;
parameter CHAN_BOND_SEQ_2_2_B = 11'b00000000000;
parameter CHAN_BOND_SEQ_2_3_A = 11'b00000000000;
parameter CHAN_BOND_SEQ_2_3_B = 11'b00000000000;
parameter CHAN_BOND_SEQ_2_4_A = 11'b00000000000;
parameter CHAN_BOND_SEQ_2_4_B = 11'b00000000000;
parameter CHAN_BOND_SEQ_2_MASK_A = 4'b1110;
parameter CHAN_BOND_SEQ_2_MASK_B = 4'b1110;
parameter CHAN_BOND_SEQ_2_USE_A = "FALSE";
parameter CHAN_BOND_SEQ_2_USE_B = "FALSE";
parameter CLK_CORRECT_USE_A = "FALSE";
parameter CLK_CORRECT_USE_B = "FALSE";
parameter CLK_COR_8B10B_DE_A = "FALSE";
parameter CLK_COR_8B10B_DE_B = "FALSE";
parameter CLK_COR_SEQ_1_1_A = 11'b00000000000;
parameter CLK_COR_SEQ_1_1_B = 11'b00000000000;
parameter CLK_COR_SEQ_1_2_A = 11'b00000000000;
parameter CLK_COR_SEQ_1_2_B = 11'b00000000000;
parameter CLK_COR_SEQ_1_3_A = 11'b00000000000;
parameter CLK_COR_SEQ_1_3_B = 11'b00000000000;
parameter CLK_COR_SEQ_1_4_A = 11'b00000000000;
parameter CLK_COR_SEQ_1_4_B = 11'b00000000000;
parameter CLK_COR_SEQ_1_MASK_A = 4'b1110;
parameter CLK_COR_SEQ_1_MASK_B = 4'b1110;
parameter CLK_COR_SEQ_2_1_A = 11'b00000000000;
parameter CLK_COR_SEQ_2_1_B = 11'b00000000000;
parameter CLK_COR_SEQ_2_2_A = 11'b00000000000;
parameter CLK_COR_SEQ_2_2_B = 11'b00000000000;
parameter CLK_COR_SEQ_2_3_A = 11'b00000000000;
parameter CLK_COR_SEQ_2_3_B = 11'b00000000000;
parameter CLK_COR_SEQ_2_4_A = 11'b00000000000;
parameter CLK_COR_SEQ_2_4_B = 11'b00000000000;
parameter CLK_COR_SEQ_2_MASK_A = 4'b1110;
parameter CLK_COR_SEQ_2_MASK_B = 4'b1110;
parameter CLK_COR_SEQ_2_USE_A = "FALSE";
parameter CLK_COR_SEQ_2_USE_B = "FALSE";
parameter CLK_COR_SEQ_DROP_A = "FALSE";
parameter CLK_COR_SEQ_DROP_B = "FALSE";
parameter COMMA32_A = "FALSE";
parameter COMMA32_B = "FALSE";
parameter COMMA_10B_MASK_A = 10'h3FF;
parameter COMMA_10B_MASK_B = 10'h3FF;
parameter CYCLE_LIMIT_SEL_A = 2'b00;
parameter CYCLE_LIMIT_SEL_B = 2'b00;
parameter DCDR_FILTER_A = 3'b010;
parameter DCDR_FILTER_B = 3'b010;
parameter DEC_MCOMMA_DETECT_A = "TRUE";
parameter DEC_MCOMMA_DETECT_B = "TRUE";
parameter DEC_PCOMMA_DETECT_A = "TRUE";
parameter DEC_PCOMMA_DETECT_B = "TRUE";
parameter DEC_VALID_COMMA_ONLY_A = "TRUE";
parameter DEC_VALID_COMMA_ONLY_B = "TRUE";
parameter DIGRX_FWDCLK_A = 2'b00;
parameter DIGRX_FWDCLK_B = 2'b00;
parameter DIGRX_SYNC_MODE_A = "FALSE";
parameter DIGRX_SYNC_MODE_B = "FALSE";
parameter ENABLE_DCDR_A = "FALSE";
parameter ENABLE_DCDR_B = "FALSE";
parameter FDET_HYS_CAL_A = 3'b010;
parameter FDET_HYS_CAL_B = 3'b010;
parameter FDET_HYS_SEL_A = 3'b100;
parameter FDET_HYS_SEL_B = 3'b100;
parameter FDET_LCK_CAL_A = 3'b100;
parameter FDET_LCK_CAL_B = 3'b100;
parameter FDET_LCK_SEL_A = 3'b001;
parameter FDET_LCK_SEL_B = 3'b001;
parameter IREFBIASMODE_A = 2'b11;
parameter IREFBIASMODE_B = 2'b11;
parameter LOOPCAL_WAIT_A = 2'b00;
parameter LOOPCAL_WAIT_B = 2'b00;
parameter MCOMMA_32B_VALUE_A = 32'h00000000;
parameter MCOMMA_32B_VALUE_B = 32'h00000000;
parameter MCOMMA_DETECT_A = "TRUE";
parameter MCOMMA_DETECT_B = "TRUE";
parameter OPPOSITE_SELECT_A = "FALSE";
parameter OPPOSITE_SELECT_B = "FALSE";
parameter PCOMMA_32B_VALUE_A = 32'h00000000;
parameter PCOMMA_32B_VALUE_B = 32'h00000000;
parameter PCOMMA_DETECT_A = "TRUE";
parameter PCOMMA_DETECT_B = "TRUE";
parameter PCS_BIT_SLIP_A = "FALSE";
parameter PCS_BIT_SLIP_B = "FALSE";
parameter PMACLKENABLE_A = "TRUE";
parameter PMACLKENABLE_B = "TRUE";
parameter PMACOREPWRENABLE_A = "TRUE";
parameter PMACOREPWRENABLE_B = "TRUE";
parameter PMAIREFTRIM_A = 4'b0111;
parameter PMAIREFTRIM_B = 4'b0111;
parameter PMAVBGCTRL_A = 5'b00000;
parameter PMAVBGCTRL_B = 5'b00000;
parameter PMAVREFTRIM_A = 4'b0111;
parameter PMAVREFTRIM_B = 4'b0111;
parameter PMA_BIT_SLIP_A = "FALSE";
parameter PMA_BIT_SLIP_B = "FALSE";
parameter POWER_ENABLE_A = "TRUE";
parameter POWER_ENABLE_B = "TRUE";
parameter REPEATER_A = "FALSE";
parameter REPEATER_B = "FALSE";
parameter RXACTST_A = "FALSE";
parameter RXACTST_B = "FALSE";
parameter RXAFEEQ_A = 9'b000000000;
parameter RXAFEEQ_B = 9'b000000000;
parameter RXAFEPD_A = "FALSE";
parameter RXAFEPD_B = "FALSE";
parameter RXAFETST_A = "FALSE";
parameter RXAFETST_B = "FALSE";
parameter RXAPD_A = "FALSE";
parameter RXAPD_B = "FALSE";
parameter RXAREGCTRL_A = 5'b00000;
parameter RXAREGCTRL_B = 5'b00000;
parameter RXASYNCDIVIDE_A = 2'b11;
parameter RXASYNCDIVIDE_B = 2'b11;
parameter RXBY_32_A = "FALSE";
parameter RXBY_32_B = "FALSE";
parameter RXCDRLOS_A = 6'b000000;
parameter RXCDRLOS_B = 6'b000000;
parameter RXCLK0_FORCE_PMACLK_A = "FALSE";
parameter RXCLK0_FORCE_PMACLK_B = "FALSE";
parameter RXCLKMODE_A = 6'b110001;
parameter RXCLKMODE_B = 6'b110001;
parameter RXCLMODE_A = 2'b00;
parameter RXCLMODE_B = 2'b00;
parameter RXCMADJ_A = 2'b01;
parameter RXCMADJ_B = 2'b01;
parameter RXCPSEL_A = "TRUE";
parameter RXCPSEL_B = "TRUE";
parameter RXCPTST_A = "FALSE";
parameter RXCPTST_B = "FALSE";
parameter RXCRCCLOCKDOUBLE_A = "FALSE";
parameter RXCRCCLOCKDOUBLE_B = "FALSE";
parameter RXCRCENABLE_A = "FALSE";
parameter RXCRCENABLE_B = "FALSE";
parameter RXCRCINITVAL_A = 32'h00000000;
parameter RXCRCINITVAL_B = 32'h00000000;
parameter RXCRCINVERTGEN_A = "FALSE";
parameter RXCRCINVERTGEN_B = "FALSE";
parameter RXCRCSAMECLOCK_A = "FALSE";
parameter RXCRCSAMECLOCK_B = "FALSE";
parameter RXCTRL1_A = 10'h200;
parameter RXCTRL1_B = 10'h200;
parameter RXCYCLE_LIMIT_SEL_A = 2'b00;
parameter RXCYCLE_LIMIT_SEL_B = 2'b00;
parameter RXDATA_SEL_A = 2'b00;
parameter RXDATA_SEL_B = 2'b00;
parameter RXDCCOUPLE_A = "FALSE";
parameter RXDCCOUPLE_B = "FALSE";
parameter RXDIGRESET_A = "FALSE";
parameter RXDIGRESET_B = "FALSE";
parameter RXDIGRX_A = "FALSE";
parameter RXDIGRX_B = "FALSE";
parameter RXEQ_A = 64'h4000000000000000;
parameter RXEQ_B = 64'h4000000000000000;
parameter RXFDCAL_CLOCK_DIVIDE_A = "NONE";
parameter RXFDCAL_CLOCK_DIVIDE_B = "NONE";
parameter RXFDET_HYS_CAL_A = 3'b010;
parameter RXFDET_HYS_CAL_B = 3'b010;
parameter RXFDET_HYS_SEL_A = 3'b100;
parameter RXFDET_HYS_SEL_B = 3'b100;
parameter RXFDET_LCK_CAL_A = 3'b100;
parameter RXFDET_LCK_CAL_B = 3'b100;
parameter RXFDET_LCK_SEL_A = 3'b001;
parameter RXFDET_LCK_SEL_B = 3'b001;
parameter RXFECONTROL1_A = 2'b00;
parameter RXFECONTROL1_B = 2'b00;
parameter RXFECONTROL2_A = 3'b000;
parameter RXFECONTROL2_B = 3'b000;
parameter RXFETUNE_A = 2'b01;
parameter RXFETUNE_B = 2'b01;
parameter RXLB_A = "FALSE";
parameter RXLB_B = "FALSE";
parameter RXLKADJ_A = 5'b00000;
parameter RXLKADJ_B = 5'b00000;
parameter RXLKAPD_A = "FALSE";
parameter RXLKAPD_B = "FALSE";
parameter RXLOOPCAL_WAIT_A = 2'b00;
parameter RXLOOPCAL_WAIT_B = 2'b00;
parameter RXLOOPFILT_A = 4'b0111;
parameter RXLOOPFILT_B = 4'b0111;
parameter RXMODE_A = 6'b000000;
parameter RXMODE_B = 6'b000000;
parameter RXPDDTST_A = "TRUE";
parameter RXPDDTST_B = "TRUE";
parameter RXPD_A = "FALSE";
parameter RXPD_B = "FALSE";
parameter RXPMACLKSEL_A = "REFCLK1";
parameter RXPMACLKSEL_B = "REFCLK1";
parameter RXRCPADJ_A = 3'b011;
parameter RXRCPADJ_B = 3'b011;
parameter RXRCPPD_A = "FALSE";
parameter RXRCPPD_B = "FALSE";
parameter RXRECCLK1_USE_SYNC_A = "FALSE";
parameter RXRECCLK1_USE_SYNC_B = "FALSE";
parameter RXRIBADJ_A = 2'b11;
parameter RXRIBADJ_B = 2'b11;
parameter RXRPDPD_A = "FALSE";
parameter RXRPDPD_B = "FALSE";
parameter RXRSDPD_A = "FALSE";
parameter RXRSDPD_B = "FALSE";
parameter RXSLOWDOWN_CAL_A = 2'b00;
parameter RXSLOWDOWN_CAL_B = 2'b00;
parameter RXTUNE_A = 13'h0000;
parameter RXTUNE_B = 13'h0000;
parameter RXVCODAC_INIT_A = 10'b1010000000;
parameter RXVCODAC_INIT_B = 10'b1010000000;
parameter RXVCO_CTRL_ENABLE_A = "FALSE";
parameter RXVCO_CTRL_ENABLE_B = "FALSE";
parameter RX_BUFFER_USE_A = "TRUE";
parameter RX_BUFFER_USE_B = "TRUE";
parameter RX_CLOCK_DIVIDER_A = 2'b00;
parameter RX_CLOCK_DIVIDER_B = 2'b00;
parameter SAMPLE_8X_A = "FALSE";
parameter SAMPLE_8X_B = "FALSE";
parameter SLOWDOWN_CAL_A = 2'b00;
parameter SLOWDOWN_CAL_B = 2'b00;
parameter TXABPMACLKSEL_A = "REFCLK1";
parameter TXABPMACLKSEL_B = "REFCLK1";
parameter TXAPD_A = "FALSE";
parameter TXAPD_B = "FALSE";
parameter TXAREFBIASSEL_A = "TRUE";
parameter TXAREFBIASSEL_B = "TRUE";
parameter TXASYNCDIVIDE_A = 2'b11;
parameter TXASYNCDIVIDE_B = 2'b11;
parameter TXCLK0_FORCE_PMACLK_A = "FALSE";
parameter TXCLK0_FORCE_PMACLK_B = "FALSE";
parameter TXCLKMODE_A = 4'b1001;
parameter TXCLKMODE_B = 4'b1001;
parameter TXCLMODE_A = 2'b00;
parameter TXCLMODE_B = 2'b00;
parameter TXCPSEL_A = "TRUE";
parameter TXCPSEL_B = "TRUE";
parameter TXCRCCLOCKDOUBLE_A = "FALSE";
parameter TXCRCCLOCKDOUBLE_B = "FALSE";
parameter TXCRCENABLE_A = "FALSE";
parameter TXCRCENABLE_B = "FALSE";
parameter TXCRCINITVAL_A = 32'h00000000;
parameter TXCRCINITVAL_B = 32'h00000000;
parameter TXCRCINVERTGEN_A = "FALSE";
parameter TXCRCINVERTGEN_B = "FALSE";
parameter TXCRCSAMECLOCK_A = "FALSE";
parameter TXCRCSAMECLOCK_B = "FALSE";
parameter TXCTRL1_A = 10'h200;
parameter TXCTRL1_B = 10'h200;
parameter TXDATA_SEL_A = 2'b00;
parameter TXDATA_SEL_B = 2'b00;
parameter TXDAT_PRDRV_DAC_A = 3'b111;
parameter TXDAT_PRDRV_DAC_B = 3'b111;
parameter TXDAT_TAP_DAC_A = 5'b10110;
parameter TXDAT_TAP_DAC_B = 5'b10110;
parameter TXDIGPD_A = "FALSE";
parameter TXDIGPD_B = "FALSE";
parameter TXFDCAL_CLOCK_DIVIDE_A = "NONE";
parameter TXFDCAL_CLOCK_DIVIDE_B = "NONE";
parameter TXHIGHSIGNALEN_A = "TRUE";
parameter TXHIGHSIGNALEN_B = "TRUE";
parameter TXLOOPFILT_A = 4'b0111;
parameter TXLOOPFILT_B = 4'b0111;
parameter TXLVLSHFTPD_A = "FALSE";
parameter TXLVLSHFTPD_B = "FALSE";
parameter TXOUTCLK1_USE_SYNC_A = "FALSE";
parameter TXOUTCLK1_USE_SYNC_B = "FALSE";
parameter TXPD_A = "FALSE";
parameter TXPD_B = "FALSE";
parameter TXPHASESEL_A = "FALSE";
parameter TXPHASESEL_B = "FALSE";
parameter TXPOST_PRDRV_DAC_A = 3'b111;
parameter TXPOST_PRDRV_DAC_B = 3'b111;
parameter TXPOST_TAP_DAC_A = 5'b01110;
parameter TXPOST_TAP_DAC_B = 5'b01110;
parameter TXPOST_TAP_PD_A = "TRUE";
parameter TXPOST_TAP_PD_B = "TRUE";
parameter TXPRE_PRDRV_DAC_A = 3'b111;
parameter TXPRE_PRDRV_DAC_B = 3'b111;
parameter TXPRE_TAP_DAC_A = 5'b00000;
parameter TXPRE_TAP_DAC_B = 5'b00000;
parameter TXPRE_TAP_PD_A = "TRUE";
parameter TXPRE_TAP_PD_B = "TRUE";
parameter TXSLEWRATE_A = "FALSE";
parameter TXSLEWRATE_B = "FALSE";
parameter TXTERMTRIM_A = 4'b1100;
parameter TXTERMTRIM_B = 4'b1100;
parameter TXTUNE_A = 13'h0000;
parameter TXTUNE_B = 13'h0000;
parameter TX_BUFFER_USE_A = "TRUE";
parameter TX_BUFFER_USE_B = "TRUE";
parameter TX_CLOCK_DIVIDER_A = 2'b00;
parameter TX_CLOCK_DIVIDER_B = 2'b00;
parameter VCODAC_INIT_A = 10'b1010000000;
parameter VCODAC_INIT_B = 10'b1010000000;
parameter VCO_CTRL_ENABLE_A = "FALSE";
parameter VCO_CTRL_ENABLE_B = "FALSE";
parameter VREFBIASMODE_A = 2'b11;
parameter VREFBIASMODE_B = 2'b11;
parameter ALIGN_COMMA_WORD_A = 4;
parameter ALIGN_COMMA_WORD_B = 4;
parameter CHAN_BOND_LIMIT_A = 16;
parameter CHAN_BOND_LIMIT_B = 16;
parameter CHAN_BOND_SEQ_LEN_A = 1;
parameter CHAN_BOND_SEQ_LEN_B = 1;
parameter CLK_COR_MAX_LAT_A = 48;
parameter CLK_COR_MAX_LAT_B = 48;
parameter CLK_COR_MIN_LAT_A = 36;
parameter CLK_COR_MIN_LAT_B = 36;
parameter CLK_COR_SEQ_LEN_A = 1;
parameter CLK_COR_SEQ_LEN_B = 1;
parameter RXOUTDIV2SEL_A = 1;
parameter RXOUTDIV2SEL_B = 1;
parameter RXPLLNDIVSEL_A = 8;
parameter RXPLLNDIVSEL_B = 8;
parameter RXUSRDIVISOR_A = 1;
parameter RXUSRDIVISOR_B = 1;
parameter SH_CNT_MAX_A = 64;
parameter SH_CNT_MAX_B = 64;
parameter SH_INVALID_CNT_MAX_A = 16;
parameter SH_INVALID_CNT_MAX_B = 16;
parameter TXOUTDIV2SEL_A = 1;
parameter TXOUTDIV2SEL_B = 1;
parameter TXPLLNDIVSEL_A = 8;
parameter TXPLLNDIVSEL_B = 8;
endmodule
//#### END MODULE DEFINITION FOR: GT11_DUAL ####

//#### BEGIN MODULE DEFINITION FOR :GTHE1_QUAD ###
module GTHE1_QUAD (
  DRDY,
  DRPDO,
  GTHINITDONE,
  MGMTPCSRDACK,
  MGMTPCSRDDATA,
  RXCODEERR0,
  RXCODEERR1,
  RXCODEERR2,
  RXCODEERR3,
  RXCTRL0,
  RXCTRL1,
  RXCTRL2,
  RXCTRL3,
  RXCTRLACK0,
  RXCTRLACK1,
  RXCTRLACK2,
  RXCTRLACK3,
  RXDATA0,
  RXDATA1,
  RXDATA2,
  RXDATA3,
  RXDATATAP0,
  RXDATATAP1,
  RXDATATAP2,
  RXDATATAP3,
  RXDISPERR0,
  RXDISPERR1,
  RXDISPERR2,
  RXDISPERR3,
  RXPCSCLKSMPL0,
  RXPCSCLKSMPL1,
  RXPCSCLKSMPL2,
  RXPCSCLKSMPL3,
  RXUSERCLKOUT0,
  RXUSERCLKOUT1,
  RXUSERCLKOUT2,
  RXUSERCLKOUT3,
  RXVALID0,
  RXVALID1,
  RXVALID2,
  RXVALID3,
  TSTPATH,
  TSTREFCLKFAB,
  TSTREFCLKOUT,
  TXCTRLACK0,
  TXCTRLACK1,
  TXCTRLACK2,
  TXCTRLACK3,
  TXDATATAP10,
  TXDATATAP11,
  TXDATATAP12,
  TXDATATAP13,
  TXDATATAP20,
  TXDATATAP21,
  TXDATATAP22,
  TXDATATAP23,
  TXN0,
  TXN1,
  TXN2,
  TXN3,
  TXP0,
  TXP1,
  TXP2,
  TXP3,
  TXPCSCLKSMPL0,
  TXPCSCLKSMPL1,
  TXPCSCLKSMPL2,
  TXPCSCLKSMPL3,
  TXUSERCLKOUT0,
  TXUSERCLKOUT1,
  TXUSERCLKOUT2,
  TXUSERCLKOUT3,
  DADDR,
  DCLK,
  DEN,
  DFETRAINCTRL0,
  DFETRAINCTRL1,
  DFETRAINCTRL2,
  DFETRAINCTRL3,
  DI,
  DISABLEDRP,
  DWE,
  GTHINIT,
  GTHRESET,
  GTHX2LANE01,
  GTHX2LANE23,
  GTHX4LANE,
  MGMTPCSLANESEL,
  MGMTPCSMMDADDR,
  MGMTPCSREGADDR,
  MGMTPCSREGRD,
  MGMTPCSREGWR,
  MGMTPCSWRDATA,
  PLLPCSCLKDIV,
  PLLREFCLKSEL,
  POWERDOWN0,
  POWERDOWN1,
  POWERDOWN2,
  POWERDOWN3,
  REFCLK,
  RXBUFRESET0,
  RXBUFRESET1,
  RXBUFRESET2,
  RXBUFRESET3,
  RXENCOMMADET0,
  RXENCOMMADET1,
  RXENCOMMADET2,
  RXENCOMMADET3,
  RXN0,
  RXN1,
  RXN2,
  RXN3,
  RXP0,
  RXP1,
  RXP2,
  RXP3,
  RXPOLARITY0,
  RXPOLARITY1,
  RXPOLARITY2,
  RXPOLARITY3,
  RXPOWERDOWN0,
  RXPOWERDOWN1,
  RXPOWERDOWN2,
  RXPOWERDOWN3,
  RXRATE0,
  RXRATE1,
  RXRATE2,
  RXRATE3,
  RXSLIP0,
  RXSLIP1,
  RXSLIP2,
  RXSLIP3,
  RXUSERCLKIN0,
  RXUSERCLKIN1,
  RXUSERCLKIN2,
  RXUSERCLKIN3,
  SAMPLERATE0,
  SAMPLERATE1,
  SAMPLERATE2,
  SAMPLERATE3,
  TXBUFRESET0,
  TXBUFRESET1,
  TXBUFRESET2,
  TXBUFRESET3,
  TXCTRL0,
  TXCTRL1,
  TXCTRL2,
  TXCTRL3,
  TXDATA0,
  TXDATA1,
  TXDATA2,
  TXDATA3,
  TXDATAMSB0,
  TXDATAMSB1,
  TXDATAMSB2,
  TXDATAMSB3,
  TXDEEMPH0,
  TXDEEMPH1,
  TXDEEMPH2,
  TXDEEMPH3,
  TXMARGIN0,
  TXMARGIN1,
  TXMARGIN2,
  TXMARGIN3,
  TXPOWERDOWN0,
  TXPOWERDOWN1,
  TXPOWERDOWN2,
  TXPOWERDOWN3,
  TXRATE0,
  TXRATE1,
  TXRATE2,
  TXRATE3,
  TXUSERCLKIN0,
  TXUSERCLKIN1,
  TXUSERCLKIN2,
  TXUSERCLKIN3
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input DCLK ;
input DEN ;
input DFETRAINCTRL0 ;
input DFETRAINCTRL1 ;
input DFETRAINCTRL2 ;
input DFETRAINCTRL3 ;
input DISABLEDRP ;
input DWE ;
input GTHINIT ;
input GTHRESET ;
input GTHX2LANE01 ;
input GTHX2LANE23 ;
input GTHX4LANE ;
input MGMTPCSREGRD ;
input MGMTPCSREGWR ;
input POWERDOWN0 ;
input POWERDOWN1 ;
input POWERDOWN2 ;
input POWERDOWN3 ;
input REFCLK ;
input RXBUFRESET0 ;
input RXBUFRESET1 ;
input RXBUFRESET2 ;
input RXBUFRESET3 ;
input RXENCOMMADET0 ;
input RXENCOMMADET1 ;
input RXENCOMMADET2 ;
input RXENCOMMADET3 ;
input RXN0 ;
input RXN1 ;
input RXN2 ;
input RXN3 ;
input RXP0 ;
input RXP1 ;
input RXP2 ;
input RXP3 ;
input RXPOLARITY0 ;
input RXPOLARITY1 ;
input RXPOLARITY2 ;
input RXPOLARITY3 ;
input RXSLIP0 ;
input RXSLIP1 ;
input RXSLIP2 ;
input RXSLIP3 ;
input RXUSERCLKIN0 ;
input RXUSERCLKIN1 ;
input RXUSERCLKIN2 ;
input RXUSERCLKIN3 ;
input TXBUFRESET0 ;
input TXBUFRESET1 ;
input TXBUFRESET2 ;
input TXBUFRESET3 ;
input TXDEEMPH0 ;
input TXDEEMPH1 ;
input TXDEEMPH2 ;
input TXDEEMPH3 ;
input TXUSERCLKIN0 ;
input TXUSERCLKIN1 ;
input TXUSERCLKIN2 ;
input TXUSERCLKIN3 ;
input [15:0] DADDR ;
input [15:0] DI ;
input [15:0] MGMTPCSREGADDR ;
input [15:0] MGMTPCSWRDATA ;
input [1:0] RXPOWERDOWN0 ;
input [1:0] RXPOWERDOWN1 ;
input [1:0] RXPOWERDOWN2 ;
input [1:0] RXPOWERDOWN3 ;
input [1:0] RXRATE0 ;
input [1:0] RXRATE1 ;
input [1:0] RXRATE2 ;
input [1:0] RXRATE3 ;
input [1:0] TXPOWERDOWN0 ;
input [1:0] TXPOWERDOWN1 ;
input [1:0] TXPOWERDOWN2 ;
input [1:0] TXPOWERDOWN3 ;
input [1:0] TXRATE0 ;
input [1:0] TXRATE1 ;
input [1:0] TXRATE2 ;
input [1:0] TXRATE3 ;
input [2:0] PLLREFCLKSEL ;
input [2:0] SAMPLERATE0 ;
input [2:0] SAMPLERATE1 ;
input [2:0] SAMPLERATE2 ;
input [2:0] SAMPLERATE3 ;
input [2:0] TXMARGIN0 ;
input [2:0] TXMARGIN1 ;
input [2:0] TXMARGIN2 ;
input [2:0] TXMARGIN3 ;
input [3:0] MGMTPCSLANESEL ;
input [4:0] MGMTPCSMMDADDR ;
input [5:0] PLLPCSCLKDIV ;
input [63:0] TXDATA0 ;
input [63:0] TXDATA1 ;
input [63:0] TXDATA2 ;
input [63:0] TXDATA3 ;
input [7:0] TXCTRL0 ;
input [7:0] TXCTRL1 ;
input [7:0] TXCTRL2 ;
input [7:0] TXCTRL3 ;
input [7:0] TXDATAMSB0 ;
input [7:0] TXDATAMSB1 ;
input [7:0] TXDATAMSB2 ;
input [7:0] TXDATAMSB3 ;
output DRDY ;
output GTHINITDONE ;
output MGMTPCSRDACK ;
output RXCTRLACK0 ;
output RXCTRLACK1 ;
output RXCTRLACK2 ;
output RXCTRLACK3 ;
output RXDATATAP0 ;
output RXDATATAP1 ;
output RXDATATAP2 ;
output RXDATATAP3 ;
output RXPCSCLKSMPL0 ;
output RXPCSCLKSMPL1 ;
output RXPCSCLKSMPL2 ;
output RXPCSCLKSMPL3 ;
output RXUSERCLKOUT0 ;
output RXUSERCLKOUT1 ;
output RXUSERCLKOUT2 ;
output RXUSERCLKOUT3 ;
output TSTPATH ;
output TSTREFCLKFAB ;
output TSTREFCLKOUT ;
output TXCTRLACK0 ;
output TXCTRLACK1 ;
output TXCTRLACK2 ;
output TXCTRLACK3 ;
output TXDATATAP10 ;
output TXDATATAP11 ;
output TXDATATAP12 ;
output TXDATATAP13 ;
output TXDATATAP20 ;
output TXDATATAP21 ;
output TXDATATAP22 ;
output TXDATATAP23 ;
output TXN0 ;
output TXN1 ;
output TXN2 ;
output TXN3 ;
output TXP0 ;
output TXP1 ;
output TXP2 ;
output TXP3 ;
output TXPCSCLKSMPL0 ;
output TXPCSCLKSMPL1 ;
output TXPCSCLKSMPL2 ;
output TXPCSCLKSMPL3 ;
output TXUSERCLKOUT0 ;
output TXUSERCLKOUT1 ;
output TXUSERCLKOUT2 ;
output TXUSERCLKOUT3 ;
output [15:0] DRPDO ;
output [15:0] MGMTPCSRDDATA ;
output [63:0] RXDATA0 ;
output [63:0] RXDATA1 ;
output [63:0] RXDATA2 ;
output [63:0] RXDATA3 ;
output [7:0] RXCODEERR0 ;
output [7:0] RXCODEERR1 ;
output [7:0] RXCODEERR2 ;
output [7:0] RXCODEERR3 ;
output [7:0] RXCTRL0 ;
output [7:0] RXCTRL1 ;
output [7:0] RXCTRL2 ;
output [7:0] RXCTRL3 ;
output [7:0] RXDISPERR0 ;
output [7:0] RXDISPERR1 ;
output [7:0] RXDISPERR2 ;
output [7:0] RXDISPERR3 ;
output [7:0] RXVALID0 ;
output [7:0] RXVALID1 ;
output [7:0] RXVALID2 ;
output [7:0] RXVALID3 ;
parameter [15:0] BER_CONST_PTRN0 = 16'h0000;
parameter [15:0] BER_CONST_PTRN1 = 16'h0000;
parameter [15:0] BUFFER_CONFIG_LANE0 = 16'h4004;
parameter [15:0] BUFFER_CONFIG_LANE1 = 16'h4004;
parameter [15:0] BUFFER_CONFIG_LANE2 = 16'h4004;
parameter [15:0] BUFFER_CONFIG_LANE3 = 16'h4004;
parameter [15:0] DFE_TRAIN_CTRL_LANE0 = 16'h0000;
parameter [15:0] DFE_TRAIN_CTRL_LANE1 = 16'h0000;
parameter [15:0] DFE_TRAIN_CTRL_LANE2 = 16'h0000;
parameter [15:0] DFE_TRAIN_CTRL_LANE3 = 16'h0000;
parameter [15:0] DLL_CFG0 = 16'h8202;
parameter [15:0] DLL_CFG1 = 16'h0000;
parameter [15:0] E10GBASEKR_LD_COEFF_UPD_LANE0 = 16'h0000;
parameter [15:0] E10GBASEKR_LD_COEFF_UPD_LANE1 = 16'h0000;
parameter [15:0] E10GBASEKR_LD_COEFF_UPD_LANE2 = 16'h0000;
parameter [15:0] E10GBASEKR_LD_COEFF_UPD_LANE3 = 16'h0000;
parameter [15:0] E10GBASEKR_LP_COEFF_UPD_LANE0 = 16'h0000;
parameter [15:0] E10GBASEKR_LP_COEFF_UPD_LANE1 = 16'h0000;
parameter [15:0] E10GBASEKR_LP_COEFF_UPD_LANE2 = 16'h0000;
parameter [15:0] E10GBASEKR_LP_COEFF_UPD_LANE3 = 16'h0000;
parameter [15:0] E10GBASEKR_PMA_CTRL_LANE0 = 16'h0002;
parameter [15:0] E10GBASEKR_PMA_CTRL_LANE1 = 16'h0002;
parameter [15:0] E10GBASEKR_PMA_CTRL_LANE2 = 16'h0002;
parameter [15:0] E10GBASEKR_PMA_CTRL_LANE3 = 16'h0002;
parameter [15:0] E10GBASEKX_CTRL_LANE0 = 16'h0000;
parameter [15:0] E10GBASEKX_CTRL_LANE1 = 16'h0000;
parameter [15:0] E10GBASEKX_CTRL_LANE2 = 16'h0000;
parameter [15:0] E10GBASEKX_CTRL_LANE3 = 16'h0000;
parameter [15:0] E10GBASER_PCS_CFG_LANE0 = 16'h070C;
parameter [15:0] E10GBASER_PCS_CFG_LANE1 = 16'h070C;
parameter [15:0] E10GBASER_PCS_CFG_LANE2 = 16'h070C;
parameter [15:0] E10GBASER_PCS_CFG_LANE3 = 16'h070C;
parameter [15:0] E10GBASER_PCS_SEEDA0_LANE0 = 16'h0001;
parameter [15:0] E10GBASER_PCS_SEEDA0_LANE1 = 16'h0001;
parameter [15:0] E10GBASER_PCS_SEEDA0_LANE2 = 16'h0001;
parameter [15:0] E10GBASER_PCS_SEEDA0_LANE3 = 16'h0001;
parameter [15:0] E10GBASER_PCS_SEEDA1_LANE0 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDA1_LANE1 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDA1_LANE2 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDA1_LANE3 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDA2_LANE0 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDA2_LANE1 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDA2_LANE2 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDA2_LANE3 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDA3_LANE0 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDA3_LANE1 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDA3_LANE2 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDA3_LANE3 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDB0_LANE0 = 16'h0001;
parameter [15:0] E10GBASER_PCS_SEEDB0_LANE1 = 16'h0001;
parameter [15:0] E10GBASER_PCS_SEEDB0_LANE2 = 16'h0001;
parameter [15:0] E10GBASER_PCS_SEEDB0_LANE3 = 16'h0001;
parameter [15:0] E10GBASER_PCS_SEEDB1_LANE0 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDB1_LANE1 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDB1_LANE2 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDB1_LANE3 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDB2_LANE0 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDB2_LANE1 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDB2_LANE2 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDB2_LANE3 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDB3_LANE0 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDB3_LANE1 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDB3_LANE2 = 16'h0000;
parameter [15:0] E10GBASER_PCS_SEEDB3_LANE3 = 16'h0000;
parameter [15:0] E10GBASER_PCS_TEST_CTRL_LANE0 = 16'h0000;
parameter [15:0] E10GBASER_PCS_TEST_CTRL_LANE1 = 16'h0000;
parameter [15:0] E10GBASER_PCS_TEST_CTRL_LANE2 = 16'h0000;
parameter [15:0] E10GBASER_PCS_TEST_CTRL_LANE3 = 16'h0000;
parameter [15:0] E10GBASEX_PCS_TSTCTRL_LANE0 = 16'h0000;
parameter [15:0] E10GBASEX_PCS_TSTCTRL_LANE1 = 16'h0000;
parameter [15:0] E10GBASEX_PCS_TSTCTRL_LANE2 = 16'h0000;
parameter [15:0] E10GBASEX_PCS_TSTCTRL_LANE3 = 16'h0000;
parameter [15:0] GLBL0_NOISE_CTRL = 16'hF0B8;
parameter [15:0] GLBL_AMON_SEL = 16'h0000;
parameter [15:0] GLBL_DMON_SEL = 16'h0200;
parameter [15:0] GLBL_PWR_CTRL = 16'h0000;
parameter [0:0] GTH_CFG_PWRUP_LANE0 = 1'b1;
parameter [0:0] GTH_CFG_PWRUP_LANE1 = 1'b1;
parameter [0:0] GTH_CFG_PWRUP_LANE2 = 1'b1;
parameter [0:0] GTH_CFG_PWRUP_LANE3 = 1'b1;
parameter [15:0] LANE_AMON_SEL = 16'h00F0;
parameter [15:0] LANE_DMON_SEL = 16'h0000;
parameter [15:0] LANE_LNK_CFGOVRD = 16'h0000;
parameter [15:0] LANE_PWR_CTRL_LANE0 = 16'h0400;
parameter [15:0] LANE_PWR_CTRL_LANE1 = 16'h0400;
parameter [15:0] LANE_PWR_CTRL_LANE2 = 16'h0400;
parameter [15:0] LANE_PWR_CTRL_LANE3 = 16'h0400;
parameter [15:0] LNK_TRN_CFG_LANE0 = 16'h0000;
parameter [15:0] LNK_TRN_CFG_LANE1 = 16'h0000;
parameter [15:0] LNK_TRN_CFG_LANE2 = 16'h0000;
parameter [15:0] LNK_TRN_CFG_LANE3 = 16'h0000;
parameter [15:0] LNK_TRN_COEFF_REQ_LANE0 = 16'h0000;
parameter [15:0] LNK_TRN_COEFF_REQ_LANE1 = 16'h0000;
parameter [15:0] LNK_TRN_COEFF_REQ_LANE2 = 16'h0000;
parameter [15:0] LNK_TRN_COEFF_REQ_LANE3 = 16'h0000;
parameter [15:0] MISC_CFG = 16'h0008;
parameter [15:0] MODE_CFG1 = 16'h0000;
parameter [15:0] MODE_CFG2 = 16'h0000;
parameter [15:0] MODE_CFG3 = 16'h0000;
parameter [15:0] MODE_CFG4 = 16'h0000;
parameter [15:0] MODE_CFG5 = 16'h0000;
parameter [15:0] MODE_CFG6 = 16'h0000;
parameter [15:0] MODE_CFG7 = 16'h0000;
parameter [15:0] PCS_ABILITY_LANE0 = 16'h0010;
parameter [15:0] PCS_ABILITY_LANE1 = 16'h0010;
parameter [15:0] PCS_ABILITY_LANE2 = 16'h0010;
parameter [15:0] PCS_ABILITY_LANE3 = 16'h0010;
parameter [15:0] PCS_CTRL1_LANE0 = 16'h2040;
parameter [15:0] PCS_CTRL1_LANE1 = 16'h2040;
parameter [15:0] PCS_CTRL1_LANE2 = 16'h2040;
parameter [15:0] PCS_CTRL1_LANE3 = 16'h2040;
parameter [15:0] PCS_CTRL2_LANE0 = 16'h0000;
parameter [15:0] PCS_CTRL2_LANE1 = 16'h0000;
parameter [15:0] PCS_CTRL2_LANE2 = 16'h0000;
parameter [15:0] PCS_CTRL2_LANE3 = 16'h0000;
parameter [15:0] PCS_MISC_CFG_0_LANE0 = 16'h1116;
parameter [15:0] PCS_MISC_CFG_0_LANE1 = 16'h1116;
parameter [15:0] PCS_MISC_CFG_0_LANE2 = 16'h1116;
parameter [15:0] PCS_MISC_CFG_0_LANE3 = 16'h1116;
parameter [15:0] PCS_MISC_CFG_1_LANE0 = 16'h0000;
parameter [15:0] PCS_MISC_CFG_1_LANE1 = 16'h0000;
parameter [15:0] PCS_MISC_CFG_1_LANE2 = 16'h0000;
parameter [15:0] PCS_MISC_CFG_1_LANE3 = 16'h0000;
parameter [15:0] PCS_MODE_LANE0 = 16'h0000;
parameter [15:0] PCS_MODE_LANE1 = 16'h0000;
parameter [15:0] PCS_MODE_LANE2 = 16'h0000;
parameter [15:0] PCS_MODE_LANE3 = 16'h0000;
parameter [15:0] PCS_RESET_1_LANE0 = 16'h0002;
parameter [15:0] PCS_RESET_1_LANE1 = 16'h0002;
parameter [15:0] PCS_RESET_1_LANE2 = 16'h0002;
parameter [15:0] PCS_RESET_1_LANE3 = 16'h0002;
parameter [15:0] PCS_RESET_LANE0 = 16'h0000;
parameter [15:0] PCS_RESET_LANE1 = 16'h0000;
parameter [15:0] PCS_RESET_LANE2 = 16'h0000;
parameter [15:0] PCS_RESET_LANE3 = 16'h0000;
parameter [15:0] PCS_TYPE_LANE0 = 16'h002C;
parameter [15:0] PCS_TYPE_LANE1 = 16'h002C;
parameter [15:0] PCS_TYPE_LANE2 = 16'h002C;
parameter [15:0] PCS_TYPE_LANE3 = 16'h002C;
parameter [15:0] PLL_CFG0 = 16'h95DF;
parameter [15:0] PLL_CFG1 = 16'h81C0;
parameter [15:0] PLL_CFG2 = 16'h0424;
parameter [15:0] PMA_CTRL1_LANE0 = 16'h0000;
parameter [15:0] PMA_CTRL1_LANE1 = 16'h0000;
parameter [15:0] PMA_CTRL1_LANE2 = 16'h0000;
parameter [15:0] PMA_CTRL1_LANE3 = 16'h0000;
parameter [15:0] PMA_CTRL2_LANE0 = 16'h000B;
parameter [15:0] PMA_CTRL2_LANE1 = 16'h000B;
parameter [15:0] PMA_CTRL2_LANE2 = 16'h000B;
parameter [15:0] PMA_CTRL2_LANE3 = 16'h000B;
parameter [15:0] PMA_LPBK_CTRL_LANE0 = 16'h0004;
parameter [15:0] PMA_LPBK_CTRL_LANE1 = 16'h0004;
parameter [15:0] PMA_LPBK_CTRL_LANE2 = 16'h0004;
parameter [15:0] PMA_LPBK_CTRL_LANE3 = 16'h0004;
parameter [15:0] PRBS_BER_CFG0_LANE0 = 16'h0000;
parameter [15:0] PRBS_BER_CFG0_LANE1 = 16'h0000;
parameter [15:0] PRBS_BER_CFG0_LANE2 = 16'h0000;
parameter [15:0] PRBS_BER_CFG0_LANE3 = 16'h0000;
parameter [15:0] PRBS_BER_CFG1_LANE0 = 16'h0000;
parameter [15:0] PRBS_BER_CFG1_LANE1 = 16'h0000;
parameter [15:0] PRBS_BER_CFG1_LANE2 = 16'h0000;
parameter [15:0] PRBS_BER_CFG1_LANE3 = 16'h0000;
parameter [15:0] PRBS_CFG_LANE0 = 16'h000A;
parameter [15:0] PRBS_CFG_LANE1 = 16'h000A;
parameter [15:0] PRBS_CFG_LANE2 = 16'h000A;
parameter [15:0] PRBS_CFG_LANE3 = 16'h000A;
parameter [15:0] PTRN_CFG0_LSB = 16'h5555;
parameter [15:0] PTRN_CFG0_MSB = 16'h5555;
parameter [15:0] PTRN_LEN_CFG = 16'h001F;
parameter [15:0] PWRUP_DLY = 16'h0000;
parameter [15:0] RX_AEQ_VAL0_LANE0 = 16'h03C0;
parameter [15:0] RX_AEQ_VAL0_LANE1 = 16'h03C0;
parameter [15:0] RX_AEQ_VAL0_LANE2 = 16'h03C0;
parameter [15:0] RX_AEQ_VAL0_LANE3 = 16'h03C0;
parameter [15:0] RX_AEQ_VAL1_LANE0 = 16'h0000;
parameter [15:0] RX_AEQ_VAL1_LANE1 = 16'h0000;
parameter [15:0] RX_AEQ_VAL1_LANE2 = 16'h0000;
parameter [15:0] RX_AEQ_VAL1_LANE3 = 16'h0000;
parameter [15:0] RX_AGC_CTRL_LANE0 = 16'h0000;
parameter [15:0] RX_AGC_CTRL_LANE1 = 16'h0000;
parameter [15:0] RX_AGC_CTRL_LANE2 = 16'h0000;
parameter [15:0] RX_AGC_CTRL_LANE3 = 16'h0000;
parameter [15:0] RX_CDR_CTRL0_LANE0 = 16'h0005;
parameter [15:0] RX_CDR_CTRL0_LANE1 = 16'h0005;
parameter [15:0] RX_CDR_CTRL0_LANE2 = 16'h0005;
parameter [15:0] RX_CDR_CTRL0_LANE3 = 16'h0005;
parameter [15:0] RX_CDR_CTRL1_LANE0 = 16'h4200;
parameter [15:0] RX_CDR_CTRL1_LANE1 = 16'h4200;
parameter [15:0] RX_CDR_CTRL1_LANE2 = 16'h4200;
parameter [15:0] RX_CDR_CTRL1_LANE3 = 16'h4200;
parameter [15:0] RX_CDR_CTRL2_LANE0 = 16'h2000;
parameter [15:0] RX_CDR_CTRL2_LANE1 = 16'h2000;
parameter [15:0] RX_CDR_CTRL2_LANE2 = 16'h2000;
parameter [15:0] RX_CDR_CTRL2_LANE3 = 16'h2000;
parameter [15:0] RX_CFG0_LANE0 = 16'h0500;
parameter [15:0] RX_CFG0_LANE1 = 16'h0500;
parameter [15:0] RX_CFG0_LANE2 = 16'h0500;
parameter [15:0] RX_CFG0_LANE3 = 16'h0500;
parameter [15:0] RX_CFG1_LANE0 = 16'h821F;
parameter [15:0] RX_CFG1_LANE1 = 16'h821F;
parameter [15:0] RX_CFG1_LANE2 = 16'h821F;
parameter [15:0] RX_CFG1_LANE3 = 16'h821F;
parameter [15:0] RX_CFG2_LANE0 = 16'h1001;
parameter [15:0] RX_CFG2_LANE1 = 16'h1001;
parameter [15:0] RX_CFG2_LANE2 = 16'h1001;
parameter [15:0] RX_CFG2_LANE3 = 16'h1001;
parameter [15:0] RX_CTLE_CTRL_LANE0 = 16'h008F;
parameter [15:0] RX_CTLE_CTRL_LANE1 = 16'h008F;
parameter [15:0] RX_CTLE_CTRL_LANE2 = 16'h008F;
parameter [15:0] RX_CTLE_CTRL_LANE3 = 16'h008F;
parameter [15:0] RX_CTRL_OVRD_LANE0 = 16'h000C;
parameter [15:0] RX_CTRL_OVRD_LANE1 = 16'h000C;
parameter [15:0] RX_CTRL_OVRD_LANE2 = 16'h000C;
parameter [15:0] RX_CTRL_OVRD_LANE3 = 16'h000C;
parameter RX_FABRIC_WIDTH0 = 6466;
parameter RX_FABRIC_WIDTH1 = 6466;
parameter RX_FABRIC_WIDTH2 = 6466;
parameter RX_FABRIC_WIDTH3 = 6466;
parameter [15:0] RX_LOOP_CTRL_LANE0 = 16'h007F;
parameter [15:0] RX_LOOP_CTRL_LANE1 = 16'h007F;
parameter [15:0] RX_LOOP_CTRL_LANE2 = 16'h007F;
parameter [15:0] RX_LOOP_CTRL_LANE3 = 16'h007F;
parameter [15:0] RX_MVAL0_LANE0 = 16'h0000;
parameter [15:0] RX_MVAL0_LANE1 = 16'h0000;
parameter [15:0] RX_MVAL0_LANE2 = 16'h0000;
parameter [15:0] RX_MVAL0_LANE3 = 16'h0000;
parameter [15:0] RX_MVAL1_LANE0 = 16'h0000;
parameter [15:0] RX_MVAL1_LANE1 = 16'h0000;
parameter [15:0] RX_MVAL1_LANE2 = 16'h0000;
parameter [15:0] RX_MVAL1_LANE3 = 16'h0000;
parameter [15:0] RX_P0S_CTRL = 16'h1206;
parameter [15:0] RX_P0_CTRL = 16'h11F0;
parameter [15:0] RX_P1_CTRL = 16'h120F;
parameter [15:0] RX_P2_CTRL = 16'h0E0F;
parameter [15:0] RX_PI_CTRL0 = 16'hD2F0;
parameter [15:0] RX_PI_CTRL1 = 16'h0080;
parameter SIM_GTHRESET_SPEEDUP = 1;
parameter SIM_VERSION = "1.0";
parameter [15:0] SLICE_CFG = 16'h0000;
parameter [15:0] SLICE_NOISE_CTRL_0_LANE01 = 16'h0000;
parameter [15:0] SLICE_NOISE_CTRL_0_LANE23 = 16'h0000;
parameter [15:0] SLICE_NOISE_CTRL_1_LANE01 = 16'h0000;
parameter [15:0] SLICE_NOISE_CTRL_1_LANE23 = 16'h0000;
parameter [15:0] SLICE_NOISE_CTRL_2_LANE01 = 16'h7FFF;
parameter [15:0] SLICE_NOISE_CTRL_2_LANE23 = 16'h7FFF;
parameter [15:0] SLICE_TX_RESET_LANE01 = 16'h0000;
parameter [15:0] SLICE_TX_RESET_LANE23 = 16'h0000;
parameter [15:0] TERM_CTRL_LANE0 = 16'h5007;
parameter [15:0] TERM_CTRL_LANE1 = 16'h5007;
parameter [15:0] TERM_CTRL_LANE2 = 16'h5007;
parameter [15:0] TERM_CTRL_LANE3 = 16'h5007;
parameter [15:0] TX_CFG0_LANE0 = 16'h203D;
parameter [15:0] TX_CFG0_LANE1 = 16'h203D;
parameter [15:0] TX_CFG0_LANE2 = 16'h203D;
parameter [15:0] TX_CFG0_LANE3 = 16'h203D;
parameter [15:0] TX_CFG1_LANE0 = 16'h0F00;
parameter [15:0] TX_CFG1_LANE1 = 16'h0F00;
parameter [15:0] TX_CFG1_LANE2 = 16'h0F00;
parameter [15:0] TX_CFG1_LANE3 = 16'h0F00;
parameter [15:0] TX_CFG2_LANE0 = 16'h0081;
parameter [15:0] TX_CFG2_LANE1 = 16'h0081;
parameter [15:0] TX_CFG2_LANE2 = 16'h0081;
parameter [15:0] TX_CFG2_LANE3 = 16'h0081;
parameter [15:0] TX_CLK_SEL0_LANE0 = 16'h2121;
parameter [15:0] TX_CLK_SEL0_LANE1 = 16'h2121;
parameter [15:0] TX_CLK_SEL0_LANE2 = 16'h2121;
parameter [15:0] TX_CLK_SEL0_LANE3 = 16'h2121;
parameter [15:0] TX_CLK_SEL1_LANE0 = 16'h2121;
parameter [15:0] TX_CLK_SEL1_LANE1 = 16'h2121;
parameter [15:0] TX_CLK_SEL1_LANE2 = 16'h2121;
parameter [15:0] TX_CLK_SEL1_LANE3 = 16'h2121;
parameter [15:0] TX_DISABLE_LANE0 = 16'h0000;
parameter [15:0] TX_DISABLE_LANE1 = 16'h0000;
parameter [15:0] TX_DISABLE_LANE2 = 16'h0000;
parameter [15:0] TX_DISABLE_LANE3 = 16'h0000;
parameter TX_FABRIC_WIDTH0 = 6466;
parameter TX_FABRIC_WIDTH1 = 6466;
parameter TX_FABRIC_WIDTH2 = 6466;
parameter TX_FABRIC_WIDTH3 = 6466;
parameter [15:0] TX_P0P0S_CTRL = 16'h060C;
parameter [15:0] TX_P1P2_CTRL = 16'h0C39;
parameter [15:0] TX_PREEMPH_LANE0 = 16'h00A1;
parameter [15:0] TX_PREEMPH_LANE1 = 16'h00A1;
parameter [15:0] TX_PREEMPH_LANE2 = 16'h00A1;
parameter [15:0] TX_PREEMPH_LANE3 = 16'h00A1;
parameter [15:0] TX_PWR_RATE_OVRD_LANE0 = 16'h0060;
parameter [15:0] TX_PWR_RATE_OVRD_LANE1 = 16'h0060;
parameter [15:0] TX_PWR_RATE_OVRD_LANE2 = 16'h0060;
parameter [15:0] TX_PWR_RATE_OVRD_LANE3 = 16'h0060;
endmodule
//#### END MODULE DEFINITION FOR: GTHE1_QUAD ####

//#### BEGIN MODULE DEFINITION FOR :GTHE2_CHANNEL ###
module GTHE2_CHANNEL (
  CPLLFBCLKLOST,
  CPLLLOCK,
  CPLLREFCLKLOST,
  DMONITOROUT,
  DRPDO,
  DRPRDY,
  EYESCANDATAERROR,
  GTHTXN,
  GTHTXP,
  GTREFCLKMONITOR,
  PCSRSVDOUT,
  PHYSTATUS,
  RSOSINTDONE,
  RXBUFSTATUS,
  RXBYTEISALIGNED,
  RXBYTEREALIGN,
  RXCDRLOCK,
  RXCHANBONDSEQ,
  RXCHANISALIGNED,
  RXCHANREALIGN,
  RXCHARISCOMMA,
  RXCHARISK,
  RXCHBONDO,
  RXCLKCORCNT,
  RXCOMINITDET,
  RXCOMMADET,
  RXCOMSASDET,
  RXCOMWAKEDET,
  RXDATA,
  RXDATAVALID,
  RXDFESLIDETAPSTARTED,
  RXDFESLIDETAPSTROBEDONE,
  RXDFESLIDETAPSTROBESTARTED,
  RXDFESTADAPTDONE,
  RXDISPERR,
  RXDLYSRESETDONE,
  RXELECIDLE,
  RXHEADER,
  RXHEADERVALID,
  RXMONITOROUT,
  RXNOTINTABLE,
  RXOSINTSTARTED,
  RXOSINTSTROBEDONE,
  RXOSINTSTROBESTARTED,
  RXOUTCLK,
  RXOUTCLKFABRIC,
  RXOUTCLKPCS,
  RXPHALIGNDONE,
  RXPHMONITOR,
  RXPHSLIPMONITOR,
  RXPMARESETDONE,
  RXPRBSERR,
  RXQPISENN,
  RXQPISENP,
  RXRATEDONE,
  RXRESETDONE,
  RXSTARTOFSEQ,
  RXSTATUS,
  RXSYNCDONE,
  RXSYNCOUT,
  RXVALID,
  TXBUFSTATUS,
  TXCOMFINISH,
  TXDLYSRESETDONE,
  TXGEARBOXREADY,
  TXOUTCLK,
  TXOUTCLKFABRIC,
  TXOUTCLKPCS,
  TXPHALIGNDONE,
  TXPHINITDONE,
  TXPMARESETDONE,
  TXQPISENN,
  TXQPISENP,
  TXRATEDONE,
  TXRESETDONE,
  TXSYNCDONE,
  TXSYNCOUT,

  CFGRESET,
  CLKRSVD0,
  CLKRSVD1,
  CPLLLOCKDETCLK,
  CPLLLOCKEN,
  CPLLPD,
  CPLLREFCLKSEL,
  CPLLRESET,
  DMONFIFORESET,
  DMONITORCLK,
  DRPADDR,
  DRPCLK,
  DRPDI,
  DRPEN,
  DRPWE,
  EYESCANMODE,
  EYESCANRESET,
  EYESCANTRIGGER,
  GTGREFCLK,
  GTHRXN,
  GTHRXP,
  GTNORTHREFCLK0,
  GTNORTHREFCLK1,
  GTREFCLK0,
  GTREFCLK1,
  GTRESETSEL,
  GTRSVD,
  GTRXRESET,
  GTSOUTHREFCLK0,
  GTSOUTHREFCLK1,
  GTTXRESET,
  LOOPBACK,
  PCSRSVDIN,
  PCSRSVDIN2,
  PMARSVDIN,
  QPLLCLK,
  QPLLREFCLK,
  RESETOVRD,
  RX8B10BEN,
  RXADAPTSELTEST,
  RXBUFRESET,
  RXCDRFREQRESET,
  RXCDRHOLD,
  RXCDROVRDEN,
  RXCDRRESET,
  RXCDRRESETRSV,
  RXCHBONDEN,
  RXCHBONDI,
  RXCHBONDLEVEL,
  RXCHBONDMASTER,
  RXCHBONDSLAVE,
  RXCOMMADETEN,
  RXDDIEN,
  RXDFEAGCHOLD,
  RXDFEAGCOVRDEN,
  RXDFEAGCTRL,
  RXDFECM1EN,
  RXDFELFHOLD,
  RXDFELFOVRDEN,
  RXDFELPMRESET,
  RXDFESLIDETAP,
  RXDFESLIDETAPADAPTEN,
  RXDFESLIDETAPHOLD,
  RXDFESLIDETAPID,
  RXDFESLIDETAPINITOVRDEN,
  RXDFESLIDETAPONLYADAPTEN,
  RXDFESLIDETAPOVRDEN,
  RXDFESLIDETAPSTROBE,
  RXDFETAP2HOLD,
  RXDFETAP2OVRDEN,
  RXDFETAP3HOLD,
  RXDFETAP3OVRDEN,
  RXDFETAP4HOLD,
  RXDFETAP4OVRDEN,
  RXDFETAP5HOLD,
  RXDFETAP5OVRDEN,
  RXDFETAP6HOLD,
  RXDFETAP6OVRDEN,
  RXDFETAP7HOLD,
  RXDFETAP7OVRDEN,
  RXDFEUTHOLD,
  RXDFEUTOVRDEN,
  RXDFEVPHOLD,
  RXDFEVPOVRDEN,
  RXDFEVSEN,
  RXDFEXYDEN,
  RXDLYBYPASS,
  RXDLYEN,
  RXDLYOVRDEN,
  RXDLYSRESET,
  RXELECIDLEMODE,
  RXGEARBOXSLIP,
  RXLPMEN,
  RXLPMHFHOLD,
  RXLPMHFOVRDEN,
  RXLPMLFHOLD,
  RXLPMLFKLOVRDEN,
  RXMCOMMAALIGNEN,
  RXMONITORSEL,
  RXOOBRESET,
  RXOSCALRESET,
  RXOSHOLD,
  RXOSINTCFG,
  RXOSINTEN,
  RXOSINTHOLD,
  RXOSINTID0,
  RXOSINTNTRLEN,
  RXOSINTOVRDEN,
  RXOSINTSTROBE,
  RXOSINTTESTOVRDEN,
  RXOSOVRDEN,
  RXOUTCLKSEL,
  RXPCOMMAALIGNEN,
  RXPCSRESET,
  RXPD,
  RXPHALIGN,
  RXPHALIGNEN,
  RXPHDLYPD,
  RXPHDLYRESET,
  RXPHOVRDEN,
  RXPMARESET,
  RXPOLARITY,
  RXPRBSCNTRESET,
  RXPRBSSEL,
  RXQPIEN,
  RXRATE,
  RXRATEMODE,
  RXSLIDE,
  RXSYNCALLIN,
  RXSYNCIN,
  RXSYNCMODE,
  RXSYSCLKSEL,
  RXUSERRDY,
  RXUSRCLK,
  RXUSRCLK2,
  SETERRSTATUS,
  SIGVALIDCLK,
  TSTIN,
  TX8B10BBYPASS,
  TX8B10BEN,
  TXBUFDIFFCTRL,
  TXCHARDISPMODE,
  TXCHARDISPVAL,
  TXCHARISK,
  TXCOMINIT,
  TXCOMSAS,
  TXCOMWAKE,
  TXDATA,
  TXDEEMPH,
  TXDETECTRX,
  TXDIFFCTRL,
  TXDIFFPD,
  TXDLYBYPASS,
  TXDLYEN,
  TXDLYHOLD,
  TXDLYOVRDEN,
  TXDLYSRESET,
  TXDLYUPDOWN,
  TXELECIDLE,
  TXHEADER,
  TXINHIBIT,
  TXMAINCURSOR,
  TXMARGIN,
  TXOUTCLKSEL,
  TXPCSRESET,
  TXPD,
  TXPDELECIDLEMODE,
  TXPHALIGN,
  TXPHALIGNEN,
  TXPHDLYPD,
  TXPHDLYRESET,
  TXPHDLYTSTCLK,
  TXPHINIT,
  TXPHOVRDEN,
  TXPIPPMEN,
  TXPIPPMOVRDEN,
  TXPIPPMPD,
  TXPIPPMSEL,
  TXPIPPMSTEPSIZE,
  TXPISOPD,
  TXPMARESET,
  TXPOLARITY,
  TXPOSTCURSOR,
  TXPOSTCURSORINV,
  TXPRBSFORCEERR,
  TXPRBSSEL,
  TXPRECURSOR,
  TXPRECURSORINV,
  TXQPIBIASEN,
  TXQPISTRONGPDOWN,
  TXQPIWEAKPUP,
  TXRATE,
  TXRATEMODE,
  TXSEQUENCE,
  TXSTARTSEQ,
  TXSWING,
  TXSYNCALLIN,
  TXSYNCIN,
  TXSYNCMODE,
  TXSYSCLKSEL,
  TXUSERRDY,
  TXUSRCLK,
  TXUSRCLK2
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CFGRESET ;
input CLKRSVD0 ;
input CLKRSVD1 ;
input CPLLLOCKDETCLK ;
input CPLLLOCKEN ;
input CPLLPD ;
input CPLLRESET ;
input DMONFIFORESET ;
input DMONITORCLK ;
input DRPCLK ;
input DRPEN ;
input DRPWE ;
input EYESCANMODE ;
input EYESCANRESET ;
input EYESCANTRIGGER ;
input GTGREFCLK ;
input GTHRXN ;
input GTHRXP ;
input GTNORTHREFCLK0 ;
input GTNORTHREFCLK1 ;
input GTREFCLK0 ;
input GTREFCLK1 ;
input GTRESETSEL ;
input GTRXRESET ;
input GTSOUTHREFCLK0 ;
input GTSOUTHREFCLK1 ;
input GTTXRESET ;
input QPLLCLK ;
input QPLLREFCLK ;
input RESETOVRD ;
input RX8B10BEN ;
input RXBUFRESET ;
input RXCDRFREQRESET ;
input RXCDRHOLD ;
input RXCDROVRDEN ;
input RXCDRRESET ;
input RXCDRRESETRSV ;
input RXCHBONDEN ;
input RXCHBONDMASTER ;
input RXCHBONDSLAVE ;
input RXCOMMADETEN ;
input RXDDIEN ;
input RXDFEAGCHOLD ;
input RXDFEAGCOVRDEN ;
input RXDFECM1EN ;
input RXDFELFHOLD ;
input RXDFELFOVRDEN ;
input RXDFELPMRESET ;
input RXDFESLIDETAPADAPTEN ;
input RXDFESLIDETAPHOLD ;
input RXDFESLIDETAPINITOVRDEN ;
input RXDFESLIDETAPONLYADAPTEN ;
input RXDFESLIDETAPOVRDEN ;
input RXDFESLIDETAPSTROBE ;
input RXDFETAP2HOLD ;
input RXDFETAP2OVRDEN ;
input RXDFETAP3HOLD ;
input RXDFETAP3OVRDEN ;
input RXDFETAP4HOLD ;
input RXDFETAP4OVRDEN ;
input RXDFETAP5HOLD ;
input RXDFETAP5OVRDEN ;
input RXDFETAP6HOLD ;
input RXDFETAP6OVRDEN ;
input RXDFETAP7HOLD ;
input RXDFETAP7OVRDEN ;
input RXDFEUTHOLD ;
input RXDFEUTOVRDEN ;
input RXDFEVPHOLD ;
input RXDFEVPOVRDEN ;
input RXDFEVSEN ;
input RXDFEXYDEN ;
input RXDLYBYPASS ;
input RXDLYEN ;
input RXDLYOVRDEN ;
input RXDLYSRESET ;
input RXGEARBOXSLIP ;
input RXLPMEN ;
input RXLPMHFHOLD ;
input RXLPMHFOVRDEN ;
input RXLPMLFHOLD ;
input RXLPMLFKLOVRDEN ;
input RXMCOMMAALIGNEN ;
input RXOOBRESET ;
input RXOSCALRESET ;
input RXOSHOLD ;
input RXOSINTEN ;
input RXOSINTHOLD ;
input RXOSINTNTRLEN ;
input RXOSINTOVRDEN ;
input RXOSINTSTROBE ;
input RXOSINTTESTOVRDEN ;
input RXOSOVRDEN ;
input RXPCOMMAALIGNEN ;
input RXPCSRESET ;
input RXPHALIGN ;
input RXPHALIGNEN ;
input RXPHDLYPD ;
input RXPHDLYRESET ;
input RXPHOVRDEN ;
input RXPMARESET ;
input RXPOLARITY ;
input RXPRBSCNTRESET ;
input RXQPIEN ;
input RXRATEMODE ;
input RXSLIDE ;
input RXSYNCALLIN ;
input RXSYNCIN ;
input RXSYNCMODE ;
input RXUSERRDY ;
input RXUSRCLK2 ;
input RXUSRCLK ;
input SETERRSTATUS ;
input SIGVALIDCLK ;
input TX8B10BEN ;
input TXCOMINIT ;
input TXCOMSAS ;
input TXCOMWAKE ;
input TXDEEMPH ;
input TXDETECTRX ;
input TXDIFFPD ;
input TXDLYBYPASS ;
input TXDLYEN ;
input TXDLYHOLD ;
input TXDLYOVRDEN ;
input TXDLYSRESET ;
input TXDLYUPDOWN ;
input TXELECIDLE ;
input TXINHIBIT ;
input TXPCSRESET ;
input TXPDELECIDLEMODE ;
input TXPHALIGN ;
input TXPHALIGNEN ;
input TXPHDLYPD ;
input TXPHDLYRESET ;
input TXPHDLYTSTCLK ;
input TXPHINIT ;
input TXPHOVRDEN ;
input TXPIPPMEN ;
input TXPIPPMOVRDEN ;
input TXPIPPMPD ;
input TXPIPPMSEL ;
input TXPISOPD ;
input TXPMARESET ;
input TXPOLARITY ;
input TXPOSTCURSORINV ;
input TXPRBSFORCEERR ;
input TXPRECURSORINV ;
input TXQPIBIASEN ;
input TXQPISTRONGPDOWN ;
input TXQPIWEAKPUP ;
input TXRATEMODE ;
input TXSTARTSEQ ;
input TXSWING ;
input TXSYNCALLIN ;
input TXSYNCIN ;
input TXSYNCMODE ;
input TXUSERRDY ;
input TXUSRCLK2 ;
input TXUSRCLK ;
input [13:0] RXADAPTSELTEST ;
input [15:0] DRPDI ;
input [15:0] GTRSVD ;
input [15:0] PCSRSVDIN ;
input [19:0] TSTIN ;
input [1:0] RXELECIDLEMODE ;
input [1:0] RXMONITORSEL ;
input [1:0] RXPD ;
input [1:0] RXSYSCLKSEL ;
input [1:0] TXPD ;
input [1:0] TXSYSCLKSEL ;
input [2:0] CPLLREFCLKSEL ;
input [2:0] LOOPBACK ;
input [2:0] RXCHBONDLEVEL ;
input [2:0] RXOUTCLKSEL ;
input [2:0] RXPRBSSEL ;
input [2:0] RXRATE ;
input [2:0] TXBUFDIFFCTRL ;
input [2:0] TXHEADER ;
input [2:0] TXMARGIN ;
input [2:0] TXOUTCLKSEL ;
input [2:0] TXPRBSSEL ;
input [2:0] TXRATE ;
input [3:0] RXOSINTCFG ;
input [3:0] RXOSINTID0 ;
input [3:0] TXDIFFCTRL ;
input [4:0] PCSRSVDIN2 ;
input [4:0] PMARSVDIN ;
input [4:0] RXCHBONDI ;
input [4:0] RXDFEAGCTRL ;
input [4:0] RXDFESLIDETAP ;
input [4:0] TXPIPPMSTEPSIZE ;
input [4:0] TXPOSTCURSOR ;
input [4:0] TXPRECURSOR ;
input [5:0] RXDFESLIDETAPID ;
input [63:0] TXDATA ;
input [6:0] TXMAINCURSOR ;
input [6:0] TXSEQUENCE ;
input [7:0] TX8B10BBYPASS ;
input [7:0] TXCHARDISPMODE ;
input [7:0] TXCHARDISPVAL ;
input [7:0] TXCHARISK ;
input [8:0] DRPADDR ;
output CPLLFBCLKLOST ;
output CPLLLOCK ;
output CPLLREFCLKLOST ;
output DRPRDY ;
output EYESCANDATAERROR ;
output GTHTXN ;
output GTHTXP ;
output GTREFCLKMONITOR ;
output PHYSTATUS ;
output RSOSINTDONE ;
output RXBYTEISALIGNED ;
output RXBYTEREALIGN ;
output RXCDRLOCK ;
output RXCHANBONDSEQ ;
output RXCHANISALIGNED ;
output RXCHANREALIGN ;
output RXCOMINITDET ;
output RXCOMMADET ;
output RXCOMSASDET ;
output RXCOMWAKEDET ;
output RXDFESLIDETAPSTARTED ;
output RXDFESLIDETAPSTROBEDONE ;
output RXDFESLIDETAPSTROBESTARTED ;
output RXDFESTADAPTDONE ;
output RXDLYSRESETDONE ;
output RXELECIDLE ;
output RXOSINTSTARTED ;
output RXOSINTSTROBEDONE ;
output RXOSINTSTROBESTARTED ;
output RXOUTCLK ;
output RXOUTCLKFABRIC ;
output RXOUTCLKPCS ;
output RXPHALIGNDONE ;
output RXPMARESETDONE ;
output RXPRBSERR ;
output RXQPISENN ;
output RXQPISENP ;
output RXRATEDONE ;
output RXRESETDONE ;
output RXSYNCDONE ;
output RXSYNCOUT ;
output RXVALID ;
output TXCOMFINISH ;
output TXDLYSRESETDONE ;
output TXGEARBOXREADY ;
output TXOUTCLK ;
output TXOUTCLKFABRIC ;
output TXOUTCLKPCS ;
output TXPHALIGNDONE ;
output TXPHINITDONE ;
output TXPMARESETDONE ;
output TXQPISENN ;
output TXQPISENP ;
output TXRATEDONE ;
output TXRESETDONE ;
output TXSYNCDONE ;
output TXSYNCOUT ;
output [14:0] DMONITOROUT ;
output [15:0] DRPDO ;
output [15:0] PCSRSVDOUT ;
output [1:0] RXCLKCORCNT ;
output [1:0] RXDATAVALID ;
output [1:0] RXHEADERVALID ;
output [1:0] RXSTARTOFSEQ ;
output [1:0] TXBUFSTATUS ;
output [2:0] RXBUFSTATUS ;
output [2:0] RXSTATUS ;
output [4:0] RXCHBONDO ;
output [4:0] RXPHMONITOR ;
output [4:0] RXPHSLIPMONITOR ;
output [5:0] RXHEADER ;
output [63:0] RXDATA ;
output [6:0] RXMONITOROUT ;
output [7:0] RXCHARISCOMMA ;
output [7:0] RXCHARISK ;
output [7:0] RXDISPERR ;
output [7:0] RXNOTINTABLE ;
parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
parameter [0:0] ACJTAG_MODE = 1'b0;
parameter [0:0] ACJTAG_RESET = 1'b0;
parameter [19:0] ADAPT_CFG0 = 20'h00C10;
parameter ALIGN_COMMA_DOUBLE = "FALSE";
parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
parameter ALIGN_COMMA_WORD = 1;
parameter ALIGN_MCOMMA_DET = "TRUE";
parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
parameter ALIGN_PCOMMA_DET = "TRUE";
parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
parameter [0:0] A_RXOSCALRESET = 1'b0;
parameter CBCC_DATA_SOURCE_SEL = "DECODED";
parameter [41:0] CFOK_CFG = 42'h24800040E80;
parameter [5:0] CFOK_CFG2 = 6'b100000;
parameter [5:0] CFOK_CFG3 = 6'b100000;
parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
parameter CHAN_BOND_MAX_SKEW = 7;
parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
parameter CHAN_BOND_SEQ_2_USE = "FALSE";
parameter CHAN_BOND_SEQ_LEN = 1;
parameter CLK_CORRECT_USE = "TRUE";
parameter CLK_COR_KEEP_IDLE = "FALSE";
parameter CLK_COR_MAX_LAT = 20;
parameter CLK_COR_MIN_LAT = 18;
parameter CLK_COR_PRECEDENCE = "TRUE";
parameter CLK_COR_REPEAT_WAIT = 0;
parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
parameter CLK_COR_SEQ_2_USE = "FALSE";
parameter CLK_COR_SEQ_LEN = 1;
parameter [28:0] CPLL_CFG = 29'h00BC07DC;
parameter CPLL_FBDIV = 4;
parameter CPLL_FBDIV_45 = 5;
parameter [23:0] CPLL_INIT_CFG = 24'h00001E;
parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
parameter CPLL_REFCLK_DIV = 1;
parameter DEC_MCOMMA_DETECT = "TRUE";
parameter DEC_PCOMMA_DETECT = "TRUE";
parameter DEC_VALID_COMMA_ONLY = "TRUE";
parameter [23:0] DMONITOR_CFG = 24'h000A00;
parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
parameter [5:0] ES_CONTROL = 6'b000000;
parameter ES_ERRDET_EN = "FALSE";
parameter ES_EYE_SCAN_EN = "TRUE";
parameter [11:0] ES_HORZ_OFFSET = 12'h000;
parameter [9:0] ES_PMA_CFG = 10'b0000000000;
parameter [4:0] ES_PRESCALE = 5'b00000;
parameter [79:0] ES_QUALIFIER = 80'h00000000000000000000;
parameter [79:0] ES_QUAL_MASK = 80'h00000000000000000000;
parameter [79:0] ES_SDATA_MASK = 80'h00000000000000000000;
parameter [8:0] ES_VERT_OFFSET = 9'b000000000;
parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
parameter FTS_LANE_DESKEW_EN = "FALSE";
parameter [2:0] GEARBOX_MODE = 3'b000;
parameter [0:0] LOOPBACK_CFG = 1'b0;
parameter [1:0] OUTREFCLK_SEL_INV = 2'b11;
parameter PCS_PCIE_EN = "FALSE";
parameter [47:0] PCS_RSVD_ATTR = 48'h000000000000;
parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
parameter [31:0] PMA_RSV = 32'b00000000000000000000000010000000;
parameter [31:0] PMA_RSV2 = 32'b00011100000000000000000000001010;
parameter [1:0] PMA_RSV3 = 2'b00;
parameter [14:0] PMA_RSV4 = 15'b000000000001000;
parameter [3:0] PMA_RSV5 = 4'b0000;
parameter [0:0] RESET_POWERSAVE_DISABLE = 1'b0;
parameter [4:0] RXBUFRESET_TIME = 5'b00001;
parameter RXBUF_ADDR_MODE = "FULL";
parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
parameter RXBUF_EN = "TRUE";
parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
parameter RXBUF_RESET_ON_EIDLE = "FALSE";
parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
parameter RXBUF_THRESH_OVFLW = 61;
parameter RXBUF_THRESH_OVRD = "FALSE";
parameter RXBUF_THRESH_UNDFLW = 4;
parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
parameter [82:0] RXCDR_CFG = 83'h0002007FE2000C208001A;
parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
parameter [5:0] RXCDR_LOCK_CFG = 6'b001001;
parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
parameter [15:0] RXDLY_CFG = 16'h001F;
parameter [8:0] RXDLY_LCFG = 9'h030;
parameter [15:0] RXDLY_TAP_CFG = 16'h0000;
parameter RXGEARBOX_EN = "FALSE";
parameter [4:0] RXISCANRESET_TIME = 5'b00001;
parameter [13:0] RXLPM_HF_CFG = 14'b00001000000000;
parameter [17:0] RXLPM_LF_CFG = 18'b001001000000000000;
parameter [6:0] RXOOB_CFG = 7'b0000110;
parameter RXOOB_CLK_CFG = "PMA";
parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
parameter [4:0] RXOSCALRESET_TIMEOUT = 5'b00000;
parameter RXOUT_DIV = 2;
parameter [4:0] RXPCSRESET_TIME = 5'b00001;
parameter [23:0] RXPHDLY_CFG = 24'h084020;
parameter [23:0] RXPH_CFG = 24'hC00002;
parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
parameter [1:0] RXPI_CFG0 = 2'b00;
parameter [1:0] RXPI_CFG1 = 2'b00;
parameter [1:0] RXPI_CFG2 = 2'b00;
parameter [1:0] RXPI_CFG3 = 2'b00;
parameter [0:0] RXPI_CFG4 = 1'b0;
parameter [0:0] RXPI_CFG5 = 1'b0;
parameter [2:0] RXPI_CFG6 = 3'b100;
parameter [4:0] RXPMARESET_TIME = 5'b00011;
parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
parameter RXSLIDE_AUTO_WAIT = 7;
parameter RXSLIDE_MODE = "OFF";
parameter [0:0] RXSYNC_MULTILANE = 1'b0;
parameter [0:0] RXSYNC_OVRD = 1'b0;
parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
parameter [23:0] RX_BIAS_CFG = 24'b000011000000000000010000;
parameter [5:0] RX_BUFFER_CFG = 6'b000000;
parameter RX_CLK25_DIV = 7;
parameter [0:0] RX_CLKMUX_PD = 1'b1;
parameter [1:0] RX_CM_SEL = 2'b11;
parameter [3:0] RX_CM_TRIM = 4'b0100;
parameter RX_DATA_WIDTH = 20;
parameter [5:0] RX_DDI_SEL = 6'b000000;
parameter [13:0] RX_DEBUG_CFG = 14'b00000000000000;
parameter RX_DEFER_RESET_BUF_EN = "TRUE";
parameter [3:0] RX_DFELPM_CFG0 = 4'b0110;
parameter [0:0] RX_DFELPM_CFG1 = 1'b0;
parameter [0:0] RX_DFELPM_KLKH_AGC_STUP_EN = 1'b1;
parameter [1:0] RX_DFE_AGC_CFG0 = 2'b00;
parameter [2:0] RX_DFE_AGC_CFG1 = 3'b010;
parameter [3:0] RX_DFE_AGC_CFG2 = 4'b0000;
parameter [0:0] RX_DFE_AGC_OVRDEN = 1'b1;
parameter [22:0] RX_DFE_GAIN_CFG = 23'h0020C0;
parameter [11:0] RX_DFE_H2_CFG = 12'b000000000000;
parameter [11:0] RX_DFE_H3_CFG = 12'b000001000000;
parameter [10:0] RX_DFE_H4_CFG = 11'b00011100000;
parameter [10:0] RX_DFE_H5_CFG = 11'b00011100000;
parameter [10:0] RX_DFE_H6_CFG = 11'b00000100000;
parameter [10:0] RX_DFE_H7_CFG = 11'b00000100000;
parameter [32:0] RX_DFE_KL_CFG = 33'b000000000000000000000001100010000;
parameter [1:0] RX_DFE_KL_LPM_KH_CFG0 = 2'b01;
parameter [2:0] RX_DFE_KL_LPM_KH_CFG1 = 3'b010;
parameter [3:0] RX_DFE_KL_LPM_KH_CFG2 = 4'b0010;
parameter [0:0] RX_DFE_KL_LPM_KH_OVRDEN = 1'b1;
parameter [1:0] RX_DFE_KL_LPM_KL_CFG0 = 2'b10;
parameter [2:0] RX_DFE_KL_LPM_KL_CFG1 = 3'b010;
parameter [3:0] RX_DFE_KL_LPM_KL_CFG2 = 4'b0010;
parameter [0:0] RX_DFE_KL_LPM_KL_OVRDEN = 1'b1;
parameter [15:0] RX_DFE_LPM_CFG = 16'h0080;
parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
parameter [53:0] RX_DFE_ST_CFG = 54'h00E100000C003F;
parameter [16:0] RX_DFE_UT_CFG = 17'b00011100000000000;
parameter [16:0] RX_DFE_VP_CFG = 17'b00011101010100011;
parameter RX_DISPERR_SEQ_MATCH = "TRUE";
parameter RX_INT_DATAWIDTH = 0;
parameter [12:0] RX_OS_CFG = 13'b0000010000000;
parameter RX_SIG_VALID_DLY = 10;
parameter RX_XCLK_SEL = "RXREC";
parameter SAS_MAX_COM = 64;
parameter SAS_MIN_COM = 36;
parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
parameter [2:0] SATA_BURST_VAL = 3'b100;
parameter SATA_CPLL_CFG = "VCO_3000MHZ";
parameter [2:0] SATA_EIDLE_VAL = 3'b100;
parameter SATA_MAX_BURST = 8;
parameter SATA_MAX_INIT = 21;
parameter SATA_MAX_WAKE = 7;
parameter SATA_MIN_BURST = 4;
parameter SATA_MIN_INIT = 12;
parameter SATA_MIN_WAKE = 4;
parameter SHOW_REALIGN_COMMA = "TRUE";
parameter [2:0] SIM_CPLLREFCLK_SEL = 3'b001;
parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
parameter SIM_RESET_SPEEDUP = "TRUE";
parameter SIM_TX_EIDLE_DRIVE_LEVEL = "X";
parameter SIM_VERSION = "1.1";
parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
parameter [2:0] TERM_RCAL_OVRD = 3'b000;
parameter [7:0] TRANS_TIME_RATE = 8'h0E;
parameter [31:0] TST_RSV = 32'h00000000;
parameter TXBUF_EN = "TRUE";
parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
parameter [15:0] TXDLY_CFG = 16'h001F;
parameter [8:0] TXDLY_LCFG = 9'h030;
parameter [15:0] TXDLY_TAP_CFG = 16'h0000;
parameter TXGEARBOX_EN = "FALSE";
parameter [0:0] TXOOB_CFG = 1'b0;
parameter TXOUT_DIV = 2;
parameter [4:0] TXPCSRESET_TIME = 5'b00001;
parameter [23:0] TXPHDLY_CFG = 24'h084020;
parameter [15:0] TXPH_CFG = 16'h0780;
parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
parameter [1:0] TXPI_CFG0 = 2'b00;
parameter [1:0] TXPI_CFG1 = 2'b00;
parameter [1:0] TXPI_CFG2 = 2'b00;
parameter [0:0] TXPI_CFG3 = 1'b0;
parameter [0:0] TXPI_CFG4 = 1'b0;
parameter [2:0] TXPI_CFG5 = 3'b100;
parameter [0:0] TXPI_GREY_SEL = 1'b0;
parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
parameter TXPI_PPMCLK_SEL = "TXUSRCLK2";
parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
parameter [4:0] TXPMARESET_TIME = 5'b00001;
parameter [0:0] TXSYNC_MULTILANE = 1'b0;
parameter [0:0] TXSYNC_OVRD = 1'b0;
parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
parameter TX_CLK25_DIV = 7;
parameter [0:0] TX_CLKMUX_PD = 1'b1;
parameter TX_DATA_WIDTH = 20;
parameter [5:0] TX_DEEMPH0 = 6'b000000;
parameter [5:0] TX_DEEMPH1 = 6'b000000;
parameter TX_DRIVE_MODE = "DIRECT";
parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
parameter TX_INT_DATAWIDTH = 0;
parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
parameter [0:0] TX_QPI_STATUS_EN = 1'b0;
parameter [13:0] TX_RXDETECT_CFG = 14'h1832;
parameter [16:0] TX_RXDETECT_PRECHARGE_TIME = 17'h00000;
parameter [2:0] TX_RXDETECT_REF = 3'b100;
parameter TX_XCLK_SEL = "TXUSR";
parameter [0:0] UCODEER_CLR = 1'b0;
parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: GTHE2_CHANNEL ####

//#### BEGIN MODULE DEFINITION FOR :GTHE2_COMMON ###
module GTHE2_COMMON (
  DRPDO,
  DRPRDY,
  PMARSVDOUT,
  QPLLDMONITOR,
  QPLLFBCLKLOST,
  QPLLLOCK,
  QPLLOUTCLK,
  QPLLOUTREFCLK,
  QPLLREFCLKLOST,
  REFCLKOUTMONITOR,

  BGBYPASSB,
  BGMONITORENB,
  BGPDB,
  BGRCALOVRD,
  BGRCALOVRDENB,
  DRPADDR,
  DRPCLK,
  DRPDI,
  DRPEN,
  DRPWE,
  GTGREFCLK,
  GTNORTHREFCLK0,
  GTNORTHREFCLK1,
  GTREFCLK0,
  GTREFCLK1,
  GTSOUTHREFCLK0,
  GTSOUTHREFCLK1,
  PMARSVD,
  QPLLLOCKDETCLK,
  QPLLLOCKEN,
  QPLLOUTRESET,
  QPLLPD,
  QPLLREFCLKSEL,
  QPLLRESET,
  QPLLRSVD1,
  QPLLRSVD2,
  RCALENB
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input BGBYPASSB ;
input BGMONITORENB ;
input BGPDB ;
input BGRCALOVRDENB ;
input DRPCLK ;
input DRPEN ;
input DRPWE ;
input GTGREFCLK ;
input GTNORTHREFCLK0 ;
input GTNORTHREFCLK1 ;
input GTREFCLK0 ;
input GTREFCLK1 ;
input GTSOUTHREFCLK0 ;
input GTSOUTHREFCLK1 ;
input QPLLLOCKDETCLK ;
input QPLLLOCKEN ;
input QPLLOUTRESET ;
input QPLLPD ;
input QPLLRESET ;
input RCALENB ;
input [15:0] DRPDI ;
input [15:0] QPLLRSVD1 ;
input [2:0] QPLLREFCLKSEL ;
input [4:0] BGRCALOVRD ;
input [4:0] QPLLRSVD2 ;
input [7:0] DRPADDR ;
input [7:0] PMARSVD ;
output DRPRDY ;
output QPLLFBCLKLOST ;
output QPLLLOCK ;
output QPLLOUTCLK ;
output QPLLOUTREFCLK ;
output QPLLREFCLKLOST ;
output REFCLKOUTMONITOR ;
output [15:0] DRPDO ;
output [15:0] PMARSVDOUT ;
output [7:0] QPLLDMONITOR ;
parameter [63:0] BIAS_CFG = 64'h0000040000001000;
parameter [31:0] COMMON_CFG = 32'h0000001C;
parameter [26:0] QPLL_CFG = 27'h0480181;
parameter [3:0] QPLL_CLKOUT_CFG = 4'b0000;
parameter [5:0] QPLL_COARSE_FREQ_OVRD = 6'b010000;
parameter [0:0] QPLL_COARSE_FREQ_OVRD_EN = 1'b0;
parameter [9:0] QPLL_CP = 10'b0000011111;
parameter [0:0] QPLL_CP_MONITOR_EN = 1'b0;
parameter [0:0] QPLL_DMONITOR_SEL = 1'b0;
parameter [9:0] QPLL_FBDIV = 10'b0000000000;
parameter [0:0] QPLL_FBDIV_MONITOR_EN = 1'b0;
parameter [0:0] QPLL_FBDIV_RATIO = 1'b0;
parameter [23:0] QPLL_INIT_CFG = 24'h000006;
parameter [15:0] QPLL_LOCK_CFG = 16'h01E8;
parameter [3:0] QPLL_LPF = 4'b1111;
parameter QPLL_REFCLK_DIV = 2;
parameter [0:0] QPLL_RP_COMP = 1'b0;
parameter [1:0] QPLL_VTRL_RESET = 2'b00;
parameter [1:0] RCAL_CFG = 2'b00;
parameter [15:0] RSVD_ATTR0 = 16'h0000;
parameter [15:0] RSVD_ATTR1 = 16'h0000;
parameter [2:0] SIM_QPLLREFCLK_SEL = 3'b001;
parameter SIM_RESET_SPEEDUP = "TRUE";
parameter SIM_VERSION = "1.1";
endmodule
//#### END MODULE DEFINITION FOR: GTHE2_COMMON ####

//#### BEGIN MODULE DEFINITION FOR :GTPA1_DUAL ###
module GTPA1_DUAL (
  DRDY,
  DRPDO,
  GTPCLKFBEAST,
  GTPCLKFBWEST,
  GTPCLKOUT0,
  GTPCLKOUT1,
  PHYSTATUS0,
  PHYSTATUS1,
  PLLLKDET0,
  PLLLKDET1,
  RCALOUTEAST,
  RCALOUTWEST,
  REFCLKOUT0,
  REFCLKOUT1,
  REFCLKPLL0,
  REFCLKPLL1,
  RESETDONE0,
  RESETDONE1,
  RXBUFSTATUS0,
  RXBUFSTATUS1,
  RXBYTEISALIGNED0,
  RXBYTEISALIGNED1,
  RXBYTEREALIGN0,
  RXBYTEREALIGN1,
  RXCHANBONDSEQ0,
  RXCHANBONDSEQ1,
  RXCHANISALIGNED0,
  RXCHANISALIGNED1,
  RXCHANREALIGN0,
  RXCHANREALIGN1,
  RXCHARISCOMMA0,
  RXCHARISCOMMA1,
  RXCHARISK0,
  RXCHARISK1,
  RXCHBONDO,
  RXCLKCORCNT0,
  RXCLKCORCNT1,
  RXCOMMADET0,
  RXCOMMADET1,
  RXDATA0,
  RXDATA1,
  RXDISPERR0,
  RXDISPERR1,
  RXELECIDLE0,
  RXELECIDLE1,
  RXLOSSOFSYNC0,
  RXLOSSOFSYNC1,
  RXNOTINTABLE0,
  RXNOTINTABLE1,
  RXPRBSERR0,
  RXPRBSERR1,
  RXRECCLK0,
  RXRECCLK1,
  RXRUNDISP0,
  RXRUNDISP1,
  RXSTATUS0,
  RXSTATUS1,
  RXVALID0,
  RXVALID1,
  TSTOUT0,
  TSTOUT1,
  TXBUFSTATUS0,
  TXBUFSTATUS1,
  TXKERR0,
  TXKERR1,
  TXN0,
  TXN1,
  TXOUTCLK0,
  TXOUTCLK1,
  TXP0,
  TXP1,
  TXRUNDISP0,
  TXRUNDISP1,
  CLK00,
  CLK01,
  CLK10,
  CLK11,
  CLKINEAST0,
  CLKINEAST1,
  CLKINWEST0,
  CLKINWEST1,
  DADDR,
  DCLK,
  DEN,
  DI,
  DWE,
  GATERXELECIDLE0,
  GATERXELECIDLE1,
  GCLK00,
  GCLK01,
  GCLK10,
  GCLK11,
  GTPCLKFBSEL0EAST,
  GTPCLKFBSEL0WEST,
  GTPCLKFBSEL1EAST,
  GTPCLKFBSEL1WEST,
  GTPRESET0,
  GTPRESET1,
  GTPTEST0,
  GTPTEST1,
  IGNORESIGDET0,
  IGNORESIGDET1,
  INTDATAWIDTH0,
  INTDATAWIDTH1,
  LOOPBACK0,
  LOOPBACK1,
  PLLCLK00,
  PLLCLK01,
  PLLCLK10,
  PLLCLK11,
  PLLLKDETEN0,
  PLLLKDETEN1,
  PLLPOWERDOWN0,
  PLLPOWERDOWN1,
  PRBSCNTRESET0,
  PRBSCNTRESET1,
  RCALINEAST,
  RCALINWEST,
  REFCLKPWRDNB0,
  REFCLKPWRDNB1,
  REFSELDYPLL0,
  REFSELDYPLL1,
  RXBUFRESET0,
  RXBUFRESET1,
  RXCDRRESET0,
  RXCDRRESET1,
  RXCHBONDI,
  RXCHBONDMASTER0,
  RXCHBONDMASTER1,
  RXCHBONDSLAVE0,
  RXCHBONDSLAVE1,
  RXCOMMADETUSE0,
  RXCOMMADETUSE1,
  RXDATAWIDTH0,
  RXDATAWIDTH1,
  RXDEC8B10BUSE0,
  RXDEC8B10BUSE1,
  RXENCHANSYNC0,
  RXENCHANSYNC1,
  RXENMCOMMAALIGN0,
  RXENMCOMMAALIGN1,
  RXENPCOMMAALIGN0,
  RXENPCOMMAALIGN1,
  RXENPMAPHASEALIGN0,
  RXENPMAPHASEALIGN1,
  RXENPRBSTST0,
  RXENPRBSTST1,
  RXEQMIX0,
  RXEQMIX1,
  RXN0,
  RXN1,
  RXP0,
  RXP1,
  RXPMASETPHASE0,
  RXPMASETPHASE1,
  RXPOLARITY0,
  RXPOLARITY1,
  RXPOWERDOWN0,
  RXPOWERDOWN1,
  RXRESET0,
  RXRESET1,
  RXSLIDE0,
  RXSLIDE1,
  RXUSRCLK0,
  RXUSRCLK1,
  RXUSRCLK20,
  RXUSRCLK21,
  TSTCLK0,
  TSTCLK1,
  TSTIN0,
  TSTIN1,
  TXBUFDIFFCTRL0,
  TXBUFDIFFCTRL1,
  TXBYPASS8B10B0,
  TXBYPASS8B10B1,
  TXCHARDISPMODE0,
  TXCHARDISPMODE1,
  TXCHARDISPVAL0,
  TXCHARDISPVAL1,
  TXCHARISK0,
  TXCHARISK1,
  TXCOMSTART0,
  TXCOMSTART1,
  TXCOMTYPE0,
  TXCOMTYPE1,
  TXDATA0,
  TXDATA1,
  TXDATAWIDTH0,
  TXDATAWIDTH1,
  TXDETECTRX0,
  TXDETECTRX1,
  TXDIFFCTRL0,
  TXDIFFCTRL1,
  TXELECIDLE0,
  TXELECIDLE1,
  TXENC8B10BUSE0,
  TXENC8B10BUSE1,
  TXENPMAPHASEALIGN0,
  TXENPMAPHASEALIGN1,
  TXENPRBSTST0,
  TXENPRBSTST1,
  TXINHIBIT0,
  TXINHIBIT1,
  TXPDOWNASYNCH0,
  TXPDOWNASYNCH1,
  TXPMASETPHASE0,
  TXPMASETPHASE1,
  TXPOLARITY0,
  TXPOLARITY1,
  TXPOWERDOWN0,
  TXPOWERDOWN1,
  TXPRBSFORCEERR0,
  TXPRBSFORCEERR1,
  TXPREEMPHASIS0,
  TXPREEMPHASIS1,
  TXRESET0,
  TXRESET1,
  TXUSRCLK0,
  TXUSRCLK1,
  TXUSRCLK20,
  TXUSRCLK21,
  USRCODEERR0,
  USRCODEERR1
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLK00 ;
input CLK01 ;
input CLK10 ;
input CLK11 ;
input CLKINEAST0 ;
input CLKINEAST1 ;
input CLKINWEST0 ;
input CLKINWEST1 ;
input DCLK ;
input DEN ;
input DWE ;
input GATERXELECIDLE0 ;
input GATERXELECIDLE1 ;
input GCLK00 ;
input GCLK01 ;
input GCLK10 ;
input GCLK11 ;
input GTPRESET0 ;
input GTPRESET1 ;
input IGNORESIGDET0 ;
input IGNORESIGDET1 ;
input INTDATAWIDTH0 ;
input INTDATAWIDTH1 ;
input PLLCLK00 ;
input PLLCLK01 ;
input PLLCLK10 ;
input PLLCLK11 ;
input PLLLKDETEN0 ;
input PLLLKDETEN1 ;
input PLLPOWERDOWN0 ;
input PLLPOWERDOWN1 ;
input PRBSCNTRESET0 ;
input PRBSCNTRESET1 ;
input REFCLKPWRDNB0 ;
input REFCLKPWRDNB1 ;
input RXBUFRESET0 ;
input RXBUFRESET1 ;
input RXCDRRESET0 ;
input RXCDRRESET1 ;
input RXCHBONDMASTER0 ;
input RXCHBONDMASTER1 ;
input RXCHBONDSLAVE0 ;
input RXCHBONDSLAVE1 ;
input RXCOMMADETUSE0 ;
input RXCOMMADETUSE1 ;
input RXDEC8B10BUSE0 ;
input RXDEC8B10BUSE1 ;
input RXENCHANSYNC0 ;
input RXENCHANSYNC1 ;
input RXENMCOMMAALIGN0 ;
input RXENMCOMMAALIGN1 ;
input RXENPCOMMAALIGN0 ;
input RXENPCOMMAALIGN1 ;
input RXENPMAPHASEALIGN0 ;
input RXENPMAPHASEALIGN1 ;
input RXN0 ;
input RXN1 ;
input RXP0 ;
input RXP1 ;
input RXPMASETPHASE0 ;
input RXPMASETPHASE1 ;
input RXPOLARITY0 ;
input RXPOLARITY1 ;
input RXRESET0 ;
input RXRESET1 ;
input RXSLIDE0 ;
input RXSLIDE1 ;
input RXUSRCLK0 ;
input RXUSRCLK1 ;
input RXUSRCLK20 ;
input RXUSRCLK21 ;
input TSTCLK0 ;
input TSTCLK1 ;
input TXCOMSTART0 ;
input TXCOMSTART1 ;
input TXCOMTYPE0 ;
input TXCOMTYPE1 ;
input TXDETECTRX0 ;
input TXDETECTRX1 ;
input TXELECIDLE0 ;
input TXELECIDLE1 ;
input TXENC8B10BUSE0 ;
input TXENC8B10BUSE1 ;
input TXENPMAPHASEALIGN0 ;
input TXENPMAPHASEALIGN1 ;
input TXINHIBIT0 ;
input TXINHIBIT1 ;
input TXPDOWNASYNCH0 ;
input TXPDOWNASYNCH1 ;
input TXPMASETPHASE0 ;
input TXPMASETPHASE1 ;
input TXPOLARITY0 ;
input TXPOLARITY1 ;
input TXPRBSFORCEERR0 ;
input TXPRBSFORCEERR1 ;
input TXRESET0 ;
input TXRESET1 ;
input TXUSRCLK0 ;
input TXUSRCLK1 ;
input TXUSRCLK20 ;
input TXUSRCLK21 ;
input USRCODEERR0 ;
input USRCODEERR1 ;
input [11:0] TSTIN0 ;
input [11:0] TSTIN1 ;
input [15:0] DI ;
input [1:0] GTPCLKFBSEL0EAST ;
input [1:0] GTPCLKFBSEL0WEST ;
input [1:0] GTPCLKFBSEL1EAST ;
input [1:0] GTPCLKFBSEL1WEST ;
input [1:0] RXDATAWIDTH0 ;
input [1:0] RXDATAWIDTH1 ;
input [1:0] RXEQMIX0 ;
input [1:0] RXEQMIX1 ;
input [1:0] RXPOWERDOWN0 ;
input [1:0] RXPOWERDOWN1 ;
input [1:0] TXDATAWIDTH0 ;
input [1:0] TXDATAWIDTH1 ;
input [1:0] TXPOWERDOWN0 ;
input [1:0] TXPOWERDOWN1 ;
input [2:0] LOOPBACK0 ;
input [2:0] LOOPBACK1 ;
input [2:0] REFSELDYPLL0 ;
input [2:0] REFSELDYPLL1 ;
input [2:0] RXCHBONDI ;
input [2:0] RXENPRBSTST0 ;
input [2:0] RXENPRBSTST1 ;
input [2:0] TXBUFDIFFCTRL0 ;
input [2:0] TXBUFDIFFCTRL1 ;
input [2:0] TXENPRBSTST0 ;
input [2:0] TXENPRBSTST1 ;
input [2:0] TXPREEMPHASIS0 ;
input [2:0] TXPREEMPHASIS1 ;
input [31:0] TXDATA0 ;
input [31:0] TXDATA1 ;
input [3:0] TXBYPASS8B10B0 ;
input [3:0] TXBYPASS8B10B1 ;
input [3:0] TXCHARDISPMODE0 ;
input [3:0] TXCHARDISPMODE1 ;
input [3:0] TXCHARDISPVAL0 ;
input [3:0] TXCHARDISPVAL1 ;
input [3:0] TXCHARISK0 ;
input [3:0] TXCHARISK1 ;
input [3:0] TXDIFFCTRL0 ;
input [3:0] TXDIFFCTRL1 ;
input [4:0] RCALINEAST ;
input [4:0] RCALINWEST ;
input [7:0] DADDR ;
input [7:0] GTPTEST0 ;
input [7:0] GTPTEST1 ;
output DRDY ;
output PHYSTATUS0 ;
output PHYSTATUS1 ;
output PLLLKDET0 ;
output PLLLKDET1 ;
output REFCLKOUT0 ;
output REFCLKOUT1 ;
output REFCLKPLL0 ;
output REFCLKPLL1 ;
output RESETDONE0 ;
output RESETDONE1 ;
output RXBYTEISALIGNED0 ;
output RXBYTEISALIGNED1 ;
output RXBYTEREALIGN0 ;
output RXBYTEREALIGN1 ;
output RXCHANBONDSEQ0 ;
output RXCHANBONDSEQ1 ;
output RXCHANISALIGNED0 ;
output RXCHANISALIGNED1 ;
output RXCHANREALIGN0 ;
output RXCHANREALIGN1 ;
output RXCOMMADET0 ;
output RXCOMMADET1 ;
output RXELECIDLE0 ;
output RXELECIDLE1 ;
output RXPRBSERR0 ;
output RXPRBSERR1 ;
output RXRECCLK0 ;
output RXRECCLK1 ;
output RXVALID0 ;
output RXVALID1 ;
output TXN0 ;
output TXN1 ;
output TXOUTCLK0 ;
output TXOUTCLK1 ;
output TXP0 ;
output TXP1 ;
output [15:0] DRPDO ;
output [1:0] GTPCLKFBEAST ;
output [1:0] GTPCLKFBWEST ;
output [1:0] GTPCLKOUT0 ;
output [1:0] GTPCLKOUT1 ;
output [1:0] RXLOSSOFSYNC0 ;
output [1:0] RXLOSSOFSYNC1 ;
output [1:0] TXBUFSTATUS0 ;
output [1:0] TXBUFSTATUS1 ;
output [2:0] RXBUFSTATUS0 ;
output [2:0] RXBUFSTATUS1 ;
output [2:0] RXCHBONDO ;
output [2:0] RXCLKCORCNT0 ;
output [2:0] RXCLKCORCNT1 ;
output [2:0] RXSTATUS0 ;
output [2:0] RXSTATUS1 ;
output [31:0] RXDATA0 ;
output [31:0] RXDATA1 ;
output [3:0] RXCHARISCOMMA0 ;
output [3:0] RXCHARISCOMMA1 ;
output [3:0] RXCHARISK0 ;
output [3:0] RXCHARISK1 ;
output [3:0] RXDISPERR0 ;
output [3:0] RXDISPERR1 ;
output [3:0] RXNOTINTABLE0 ;
output [3:0] RXNOTINTABLE1 ;
output [3:0] RXRUNDISP0 ;
output [3:0] RXRUNDISP1 ;
output [3:0] TXKERR0 ;
output [3:0] TXKERR1 ;
output [3:0] TXRUNDISP0 ;
output [3:0] TXRUNDISP1 ;
output [4:0] RCALOUTEAST ;
output [4:0] RCALOUTWEST ;
output [4:0] TSTOUT0 ;
output [4:0] TSTOUT1 ;
parameter AC_CAP_DIS_0 = "TRUE";
parameter AC_CAP_DIS_1 = "TRUE";
parameter ALIGN_COMMA_WORD_0 = 1;
parameter ALIGN_COMMA_WORD_1 = 1;
parameter CB2_INH_CC_PERIOD_0 = 8;
parameter CB2_INH_CC_PERIOD_1 = 8;
parameter [4:0] CDR_PH_ADJ_TIME_0 = 5'b01010;
parameter [4:0] CDR_PH_ADJ_TIME_1 = 5'b01010;
parameter CHAN_BOND_1_MAX_SKEW_0 = 7;
parameter CHAN_BOND_1_MAX_SKEW_1 = 7;
parameter CHAN_BOND_2_MAX_SKEW_0 = 1;
parameter CHAN_BOND_2_MAX_SKEW_1 = 1;
parameter CHAN_BOND_KEEP_ALIGN_0 = "FALSE";
parameter CHAN_BOND_KEEP_ALIGN_1 = "FALSE";
parameter [9:0] CHAN_BOND_SEQ_1_1_0 = 10'b0101111100;
parameter [9:0] CHAN_BOND_SEQ_1_1_1 = 10'b0101111100;
parameter [9:0] CHAN_BOND_SEQ_1_2_0 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_2_1 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_3_0 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_3_1 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_4_0 = 10'b0110111100;
parameter [9:0] CHAN_BOND_SEQ_1_4_1 = 10'b0110111100;
parameter [3:0] CHAN_BOND_SEQ_1_ENABLE_0 = 4'b1111;
parameter [3:0] CHAN_BOND_SEQ_1_ENABLE_1 = 4'b1111;
parameter [9:0] CHAN_BOND_SEQ_2_1_0 = 10'b0110111100;
parameter [9:0] CHAN_BOND_SEQ_2_1_1 = 10'b0110111100;
parameter [9:0] CHAN_BOND_SEQ_2_2_0 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_2_1 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_3_0 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_3_1 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_4_0 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_4_1 = 10'b0100111100;
parameter [3:0] CHAN_BOND_SEQ_2_ENABLE_0 = 4'b1111;
parameter [3:0] CHAN_BOND_SEQ_2_ENABLE_1 = 4'b1111;
parameter CHAN_BOND_SEQ_2_USE_0 = "FALSE";
parameter CHAN_BOND_SEQ_2_USE_1 = "FALSE";
parameter CHAN_BOND_SEQ_LEN_0 = 1;
parameter CHAN_BOND_SEQ_LEN_1 = 1;
parameter CLK25_DIVIDER_0 = 4;
parameter CLK25_DIVIDER_1 = 4;
parameter CLKINDC_B_0 = "TRUE";
parameter CLKINDC_B_1 = "TRUE";
parameter CLKRCV_TRST_0 = "TRUE";
parameter CLKRCV_TRST_1 = "TRUE";
parameter CLK_CORRECT_USE_0 = "TRUE";
parameter CLK_CORRECT_USE_1 = "TRUE";
parameter CLK_COR_ADJ_LEN_0 = 1;
parameter CLK_COR_ADJ_LEN_1 = 1;
parameter CLK_COR_DET_LEN_0 = 1;
parameter CLK_COR_DET_LEN_1 = 1;
parameter CLK_COR_INSERT_IDLE_FLAG_0 = "FALSE";
parameter CLK_COR_INSERT_IDLE_FLAG_1 = "FALSE";
parameter CLK_COR_KEEP_IDLE_0 = "FALSE";
parameter CLK_COR_KEEP_IDLE_1 = "FALSE";
parameter CLK_COR_MAX_LAT_0 = 20;
parameter CLK_COR_MAX_LAT_1 = 20;
parameter CLK_COR_MIN_LAT_0 = 18;
parameter CLK_COR_MIN_LAT_1 = 18;
parameter CLK_COR_PRECEDENCE_0 = "TRUE";
parameter CLK_COR_PRECEDENCE_1 = "TRUE";
parameter CLK_COR_REPEAT_WAIT_0 = 0;
parameter CLK_COR_REPEAT_WAIT_1 = 0;
parameter [9:0] CLK_COR_SEQ_1_1_0 = 10'b0100011100;
parameter [9:0] CLK_COR_SEQ_1_1_1 = 10'b0100011100;
parameter [9:0] CLK_COR_SEQ_1_2_0 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_2_1 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_3_0 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_3_1 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_4_0 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_4_1 = 10'b0000000000;
parameter [3:0] CLK_COR_SEQ_1_ENABLE_0 = 4'b1111;
parameter [3:0] CLK_COR_SEQ_1_ENABLE_1 = 4'b1111;
parameter [9:0] CLK_COR_SEQ_2_1_0 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_1_1 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_2_0 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_2_1 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_3_0 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_3_1 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_4_0 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_4_1 = 10'b0000000000;
parameter [3:0] CLK_COR_SEQ_2_ENABLE_0 = 4'b1111;
parameter [3:0] CLK_COR_SEQ_2_ENABLE_1 = 4'b1111;
parameter CLK_COR_SEQ_2_USE_0 = "FALSE";
parameter CLK_COR_SEQ_2_USE_1 = "FALSE";
parameter CLK_OUT_GTP_SEL_0 = "REFCLKPLL0";
parameter CLK_OUT_GTP_SEL_1 = "REFCLKPLL1";
parameter [1:0] CM_TRIM_0 = 2'b00;
parameter [1:0] CM_TRIM_1 = 2'b00;
parameter [9:0] COMMA_10B_ENABLE_0 = 10'b1111111111;
parameter [9:0] COMMA_10B_ENABLE_1 = 10'b1111111111;
parameter [3:0] COM_BURST_VAL_0 = 4'b1111;
parameter [3:0] COM_BURST_VAL_1 = 4'b1111;
parameter DEC_MCOMMA_DETECT_0 = "TRUE";
parameter DEC_MCOMMA_DETECT_1 = "TRUE";
parameter DEC_PCOMMA_DETECT_0 = "TRUE";
parameter DEC_PCOMMA_DETECT_1 = "TRUE";
parameter DEC_VALID_COMMA_ONLY_0 = "TRUE";
parameter DEC_VALID_COMMA_ONLY_1 = "TRUE";
parameter GTP_CFG_PWRUP_0 = "TRUE";
parameter GTP_CFG_PWRUP_1 = "TRUE";
parameter [9:0] MCOMMA_10B_VALUE_0 = 10'b1010000011;
parameter [9:0] MCOMMA_10B_VALUE_1 = 10'b1010000011;
parameter MCOMMA_DETECT_0 = "TRUE";
parameter MCOMMA_DETECT_1 = "TRUE";
parameter [2:0] OOBDETECT_THRESHOLD_0 = 3'b110;
parameter [2:0] OOBDETECT_THRESHOLD_1 = 3'b110;
parameter OOB_CLK_DIVIDER_0 = 4;
parameter OOB_CLK_DIVIDER_1 = 4;
parameter PCI_EXPRESS_MODE_0 = "FALSE";
parameter PCI_EXPRESS_MODE_1 = "FALSE";
parameter [9:0] PCOMMA_10B_VALUE_0 = 10'b0101111100;
parameter [9:0] PCOMMA_10B_VALUE_1 = 10'b0101111100;
parameter PCOMMA_DETECT_0 = "TRUE";
parameter PCOMMA_DETECT_1 = "TRUE";
parameter [2:0] PLLLKDET_CFG_0 = 3'b101;
parameter [2:0] PLLLKDET_CFG_1 = 3'b101;
parameter [23:0] PLL_COM_CFG_0 = 24'h21680A;
parameter [23:0] PLL_COM_CFG_1 = 24'h21680A;
parameter [7:0] PLL_CP_CFG_0 = 8'h00;
parameter [7:0] PLL_CP_CFG_1 = 8'h00;
parameter PLL_DIVSEL_FB_0 = 5;
parameter PLL_DIVSEL_FB_1 = 5;
parameter PLL_DIVSEL_REF_0 = 2;
parameter PLL_DIVSEL_REF_1 = 2;
parameter PLL_RXDIVSEL_OUT_0 = 1;
parameter PLL_RXDIVSEL_OUT_1 = 1;
parameter PLL_SATA_0 = "FALSE";
parameter PLL_SATA_1 = "FALSE";
parameter PLL_SOURCE_0 = "PLL0";
parameter PLL_SOURCE_1 = "PLL0";
parameter PLL_TXDIVSEL_OUT_0 = 1;
parameter PLL_TXDIVSEL_OUT_1 = 1;
parameter [26:0] PMA_CDR_SCAN_0 = 27'h6404040;
parameter [26:0] PMA_CDR_SCAN_1 = 27'h6404040;
parameter [35:0] PMA_COM_CFG_EAST = 36'h000008000;
parameter [35:0] PMA_COM_CFG_WEST = 36'h00000A000;
parameter [6:0] PMA_RXSYNC_CFG_0 = 7'h00;
parameter [6:0] PMA_RXSYNC_CFG_1 = 7'h00;
parameter [24:0] PMA_RX_CFG_0 = 25'h05CE048;
parameter [24:0] PMA_RX_CFG_1 = 25'h05CE048;
parameter [19:0] PMA_TX_CFG_0 = 20'h00082;
parameter [19:0] PMA_TX_CFG_1 = 20'h00082;
parameter RCV_TERM_GND_0 = "FALSE";
parameter RCV_TERM_GND_1 = "FALSE";
parameter RCV_TERM_VTTRX_0 = "TRUE";
parameter RCV_TERM_VTTRX_1 = "TRUE";
parameter [7:0] RXEQ_CFG_0 = 8'b01111011;
parameter [7:0] RXEQ_CFG_1 = 8'b01111011;
parameter [0:0] RXPRBSERR_LOOPBACK_0 = 1'b0;
parameter [0:0] RXPRBSERR_LOOPBACK_1 = 1'b0;
parameter RX_BUFFER_USE_0 = "TRUE";
parameter RX_BUFFER_USE_1 = "TRUE";
parameter RX_DECODE_SEQ_MATCH_0 = "TRUE";
parameter RX_DECODE_SEQ_MATCH_1 = "TRUE";
parameter RX_EN_IDLE_HOLD_CDR_0 = "FALSE";
parameter RX_EN_IDLE_HOLD_CDR_1 = "FALSE";
parameter RX_EN_IDLE_RESET_BUF_0 = "TRUE";
parameter RX_EN_IDLE_RESET_BUF_1 = "TRUE";
parameter RX_EN_IDLE_RESET_FR_0 = "TRUE";
parameter RX_EN_IDLE_RESET_FR_1 = "TRUE";
parameter RX_EN_IDLE_RESET_PH_0 = "TRUE";
parameter RX_EN_IDLE_RESET_PH_1 = "TRUE";
parameter RX_EN_MODE_RESET_BUF_0 = "TRUE";
parameter RX_EN_MODE_RESET_BUF_1 = "TRUE";
parameter [3:0] RX_IDLE_HI_CNT_0 = 4'b1000;
parameter [3:0] RX_IDLE_HI_CNT_1 = 4'b1000;
parameter [3:0] RX_IDLE_LO_CNT_0 = 4'b0000;
parameter [3:0] RX_IDLE_LO_CNT_1 = 4'b0000;
parameter RX_LOSS_OF_SYNC_FSM_0 = "FALSE";
parameter RX_LOSS_OF_SYNC_FSM_1 = "FALSE";
parameter RX_LOS_INVALID_INCR_0 = 1;
parameter RX_LOS_INVALID_INCR_1 = 1;
parameter RX_LOS_THRESHOLD_0 = 4;
parameter RX_LOS_THRESHOLD_1 = 4;
parameter RX_SLIDE_MODE_0 = "PCS";
parameter RX_SLIDE_MODE_1 = "PCS";
parameter RX_STATUS_FMT_0 = "PCIE";
parameter RX_STATUS_FMT_1 = "PCIE";
parameter RX_XCLK_SEL_0 = "RXREC";
parameter RX_XCLK_SEL_1 = "RXREC";
parameter [2:0] SATA_BURST_VAL_0 = 3'b100;
parameter [2:0] SATA_BURST_VAL_1 = 3'b100;
parameter [2:0] SATA_IDLE_VAL_0 = 3'b011;
parameter [2:0] SATA_IDLE_VAL_1 = 3'b011;
parameter SATA_MAX_BURST_0 = 7;
parameter SATA_MAX_BURST_1 = 7;
parameter SATA_MAX_INIT_0 = 22;
parameter SATA_MAX_INIT_1 = 22;
parameter SATA_MAX_WAKE_0 = 7;
parameter SATA_MAX_WAKE_1 = 7;
parameter SATA_MIN_BURST_0 = 4;
parameter SATA_MIN_BURST_1 = 4;
parameter SATA_MIN_INIT_0 = 12;
parameter SATA_MIN_INIT_1 = 12;
parameter SATA_MIN_WAKE_0 = 4;
parameter SATA_MIN_WAKE_1 = 4;
parameter SIM_GTPRESET_SPEEDUP = 0;
parameter SIM_RECEIVER_DETECT_PASS = "FALSE";
parameter [2:0] SIM_REFCLK0_SOURCE = 3'b000;
parameter [2:0] SIM_REFCLK1_SOURCE = 3'b000;
parameter SIM_TX_ELEC_IDLE_LEVEL = "X";
parameter SIM_VERSION = "2.0";
parameter [4:0] TERMINATION_CTRL_0 = 5'b10100;
parameter [4:0] TERMINATION_CTRL_1 = 5'b10100;
parameter TERMINATION_OVRD_0 = "FALSE";
parameter TERMINATION_OVRD_1 = "FALSE";
parameter [11:0] TRANS_TIME_FROM_P2_0 = 12'h03C;
parameter [11:0] TRANS_TIME_FROM_P2_1 = 12'h03C;
parameter [7:0] TRANS_TIME_NON_P2_0 = 8'h19;
parameter [7:0] TRANS_TIME_NON_P2_1 = 8'h19;
parameter [9:0] TRANS_TIME_TO_P2_0 = 10'h064;
parameter [9:0] TRANS_TIME_TO_P2_1 = 10'h064;
parameter [31:0] TST_ATTR_0 = 32'h00000000;
parameter [31:0] TST_ATTR_1 = 32'h00000000;
parameter [2:0] TXRX_INVERT_0 = 3'b011;
parameter [2:0] TXRX_INVERT_1 = 3'b011;
parameter TX_BUFFER_USE_0 = "FALSE";
parameter TX_BUFFER_USE_1 = "FALSE";
parameter [13:0] TX_DETECT_RX_CFG_0 = 14'h1832;
parameter [13:0] TX_DETECT_RX_CFG_1 = 14'h1832;
parameter [2:0] TX_IDLE_DELAY_0 = 3'b011;
parameter [2:0] TX_IDLE_DELAY_1 = 3'b011;
parameter [1:0] TX_TDCC_CFG_0 = 2'b00;
parameter [1:0] TX_TDCC_CFG_1 = 2'b00;
parameter TX_XCLK_SEL_0 = "TXUSR";
parameter TX_XCLK_SEL_1 = "TXUSR";
endmodule
//#### END MODULE DEFINITION FOR: GTPA1_DUAL ####

//#### BEGIN MODULE DEFINITION FOR :GTPE2_CHANNEL ###
module GTPE2_CHANNEL (
  DMONITOROUT,
  DRPDO,
  DRPRDY,
  EYESCANDATAERROR,
  GTPTXN,
  GTPTXP,
  PCSRSVDOUT,
  PHYSTATUS,
  PMARSVDOUT0,
  PMARSVDOUT1,
  RXBUFSTATUS,
  RXBYTEISALIGNED,
  RXBYTEREALIGN,
  RXCDRLOCK,
  RXCHANBONDSEQ,
  RXCHANISALIGNED,
  RXCHANREALIGN,
  RXCHARISCOMMA,
  RXCHARISK,
  RXCHBONDO,
  RXCLKCORCNT,
  RXCOMINITDET,
  RXCOMMADET,
  RXCOMSASDET,
  RXCOMWAKEDET,
  RXDATA,
  RXDATAVALID,
  RXDISPERR,
  RXDLYSRESETDONE,
  RXELECIDLE,
  RXHEADER,
  RXHEADERVALID,
  RXNOTINTABLE,
  RXOSINTDONE,
  RXOSINTSTARTED,
  RXOSINTSTROBEDONE,
  RXOSINTSTROBESTARTED,
  RXOUTCLK,
  RXOUTCLKFABRIC,
  RXOUTCLKPCS,
  RXPHALIGNDONE,
  RXPHMONITOR,
  RXPHSLIPMONITOR,
  RXPMARESETDONE,
  RXPRBSERR,
  RXRATEDONE,
  RXRESETDONE,
  RXSTARTOFSEQ,
  RXSTATUS,
  RXSYNCDONE,
  RXSYNCOUT,
  RXVALID,
  TXBUFSTATUS,
  TXCOMFINISH,
  TXDLYSRESETDONE,
  TXGEARBOXREADY,
  TXOUTCLK,
  TXOUTCLKFABRIC,
  TXOUTCLKPCS,
  TXPHALIGNDONE,
  TXPHINITDONE,
  TXPMARESETDONE,
  TXRATEDONE,
  TXRESETDONE,
  TXSYNCDONE,
  TXSYNCOUT,

  CFGRESET,
  CLKRSVD0,
  CLKRSVD1,
  DMONFIFORESET,
  DMONITORCLK,
  DRPADDR,
  DRPCLK,
  DRPDI,
  DRPEN,
  DRPWE,
  EYESCANMODE,
  EYESCANRESET,
  EYESCANTRIGGER,
  GTPRXN,
  GTPRXP,
  GTRESETSEL,
  GTRSVD,
  GTRXRESET,
  GTTXRESET,
  LOOPBACK,
  PCSRSVDIN,
  PLL0CLK,
  PLL0REFCLK,
  PLL1CLK,
  PLL1REFCLK,
  PMARSVDIN0,
  PMARSVDIN1,
  PMARSVDIN2,
  PMARSVDIN3,
  PMARSVDIN4,
  RESETOVRD,
  RX8B10BEN,
  RXADAPTSELTEST,
  RXBUFRESET,
  RXCDRFREQRESET,
  RXCDRHOLD,
  RXCDROVRDEN,
  RXCDRRESET,
  RXCDRRESETRSV,
  RXCHBONDEN,
  RXCHBONDI,
  RXCHBONDLEVEL,
  RXCHBONDMASTER,
  RXCHBONDSLAVE,
  RXCOMMADETEN,
  RXDDIEN,
  RXDFEXYDEN,
  RXDLYBYPASS,
  RXDLYEN,
  RXDLYOVRDEN,
  RXDLYSRESET,
  RXELECIDLEMODE,
  RXGEARBOXSLIP,
  RXLPMHFHOLD,
  RXLPMHFOVRDEN,
  RXLPMLFHOLD,
  RXLPMLFOVRDEN,
  RXLPMOSINTNTRLEN,
  RXLPMRESET,
  RXMCOMMAALIGNEN,
  RXOOBRESET,
  RXOSCALRESET,
  RXOSHOLD,
  RXOSINTCFG,
  RXOSINTEN,
  RXOSINTHOLD,
  RXOSINTID0,
  RXOSINTNTRLEN,
  RXOSINTOVRDEN,
  RXOSINTPD,
  RXOSINTSTROBE,
  RXOSINTTESTOVRDEN,
  RXOSOVRDEN,
  RXOUTCLKSEL,
  RXPCOMMAALIGNEN,
  RXPCSRESET,
  RXPD,
  RXPHALIGN,
  RXPHALIGNEN,
  RXPHDLYPD,
  RXPHDLYRESET,
  RXPHOVRDEN,
  RXPMARESET,
  RXPOLARITY,
  RXPRBSCNTRESET,
  RXPRBSSEL,
  RXRATE,
  RXRATEMODE,
  RXSLIDE,
  RXSYNCALLIN,
  RXSYNCIN,
  RXSYNCMODE,
  RXSYSCLKSEL,
  RXUSERRDY,
  RXUSRCLK,
  RXUSRCLK2,
  SETERRSTATUS,
  SIGVALIDCLK,
  TSTIN,
  TX8B10BBYPASS,
  TX8B10BEN,
  TXBUFDIFFCTRL,
  TXCHARDISPMODE,
  TXCHARDISPVAL,
  TXCHARISK,
  TXCOMINIT,
  TXCOMSAS,
  TXCOMWAKE,
  TXDATA,
  TXDEEMPH,
  TXDETECTRX,
  TXDIFFCTRL,
  TXDIFFPD,
  TXDLYBYPASS,
  TXDLYEN,
  TXDLYHOLD,
  TXDLYOVRDEN,
  TXDLYSRESET,
  TXDLYUPDOWN,
  TXELECIDLE,
  TXHEADER,
  TXINHIBIT,
  TXMAINCURSOR,
  TXMARGIN,
  TXOUTCLKSEL,
  TXPCSRESET,
  TXPD,
  TXPDELECIDLEMODE,
  TXPHALIGN,
  TXPHALIGNEN,
  TXPHDLYPD,
  TXPHDLYRESET,
  TXPHDLYTSTCLK,
  TXPHINIT,
  TXPHOVRDEN,
  TXPIPPMEN,
  TXPIPPMOVRDEN,
  TXPIPPMPD,
  TXPIPPMSEL,
  TXPIPPMSTEPSIZE,
  TXPISOPD,
  TXPMARESET,
  TXPOLARITY,
  TXPOSTCURSOR,
  TXPOSTCURSORINV,
  TXPRBSFORCEERR,
  TXPRBSSEL,
  TXPRECURSOR,
  TXPRECURSORINV,
  TXRATE,
  TXRATEMODE,
  TXSEQUENCE,
  TXSTARTSEQ,
  TXSWING,
  TXSYNCALLIN,
  TXSYNCIN,
  TXSYNCMODE,
  TXSYSCLKSEL,
  TXUSERRDY,
  TXUSRCLK,
  TXUSRCLK2
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CFGRESET ;
input CLKRSVD0 ;
input CLKRSVD1 ;
input DMONFIFORESET ;
input DMONITORCLK ;
input DRPCLK ;
input DRPEN ;
input DRPWE ;
input EYESCANMODE ;
input EYESCANRESET ;
input EYESCANTRIGGER ;
input GTPRXN ;
input GTPRXP ;
input GTRESETSEL ;
input GTRXRESET ;
input GTTXRESET ;
input PLL0CLK ;
input PLL0REFCLK ;
input PLL1CLK ;
input PLL1REFCLK ;
input PMARSVDIN0 ;
input PMARSVDIN1 ;
input PMARSVDIN2 ;
input PMARSVDIN3 ;
input PMARSVDIN4 ;
input RESETOVRD ;
input RX8B10BEN ;
input RXBUFRESET ;
input RXCDRFREQRESET ;
input RXCDRHOLD ;
input RXCDROVRDEN ;
input RXCDRRESET ;
input RXCDRRESETRSV ;
input RXCHBONDEN ;
input RXCHBONDMASTER ;
input RXCHBONDSLAVE ;
input RXCOMMADETEN ;
input RXDDIEN ;
input RXDFEXYDEN ;
input RXDLYBYPASS ;
input RXDLYEN ;
input RXDLYOVRDEN ;
input RXDLYSRESET ;
input RXGEARBOXSLIP ;
input RXLPMHFHOLD ;
input RXLPMHFOVRDEN ;
input RXLPMLFHOLD ;
input RXLPMLFOVRDEN ;
input RXLPMOSINTNTRLEN ;
input RXLPMRESET ;
input RXMCOMMAALIGNEN ;
input RXOOBRESET ;
input RXOSCALRESET ;
input RXOSHOLD ;
input RXOSINTEN ;
input RXOSINTHOLD ;
input RXOSINTNTRLEN ;
input RXOSINTOVRDEN ;
input RXOSINTPD ;
input RXOSINTSTROBE ;
input RXOSINTTESTOVRDEN ;
input RXOSOVRDEN ;
input RXPCOMMAALIGNEN ;
input RXPCSRESET ;
input RXPHALIGN ;
input RXPHALIGNEN ;
input RXPHDLYPD ;
input RXPHDLYRESET ;
input RXPHOVRDEN ;
input RXPMARESET ;
input RXPOLARITY ;
input RXPRBSCNTRESET ;
input RXRATEMODE ;
input RXSLIDE ;
input RXSYNCALLIN ;
input RXSYNCIN ;
input RXSYNCMODE ;
input RXUSERRDY ;
input RXUSRCLK2 ;
input RXUSRCLK ;
input SETERRSTATUS ;
input SIGVALIDCLK ;
input TX8B10BEN ;
input TXCOMINIT ;
input TXCOMSAS ;
input TXCOMWAKE ;
input TXDEEMPH ;
input TXDETECTRX ;
input TXDIFFPD ;
input TXDLYBYPASS ;
input TXDLYEN ;
input TXDLYHOLD ;
input TXDLYOVRDEN ;
input TXDLYSRESET ;
input TXDLYUPDOWN ;
input TXELECIDLE ;
input TXINHIBIT ;
input TXPCSRESET ;
input TXPDELECIDLEMODE ;
input TXPHALIGN ;
input TXPHALIGNEN ;
input TXPHDLYPD ;
input TXPHDLYRESET ;
input TXPHDLYTSTCLK ;
input TXPHINIT ;
input TXPHOVRDEN ;
input TXPIPPMEN ;
input TXPIPPMOVRDEN ;
input TXPIPPMPD ;
input TXPIPPMSEL ;
input TXPISOPD ;
input TXPMARESET ;
input TXPOLARITY ;
input TXPOSTCURSORINV ;
input TXPRBSFORCEERR ;
input TXPRECURSORINV ;
input TXRATEMODE ;
input TXSTARTSEQ ;
input TXSWING ;
input TXSYNCALLIN ;
input TXSYNCIN ;
input TXSYNCMODE ;
input TXUSERRDY ;
input TXUSRCLK2 ;
input TXUSRCLK ;
input [13:0] RXADAPTSELTEST ;
input [15:0] DRPDI ;
input [15:0] GTRSVD ;
input [15:0] PCSRSVDIN ;
input [19:0] TSTIN ;
input [1:0] RXELECIDLEMODE ;
input [1:0] RXPD ;
input [1:0] RXSYSCLKSEL ;
input [1:0] TXPD ;
input [1:0] TXSYSCLKSEL ;
input [2:0] LOOPBACK ;
input [2:0] RXCHBONDLEVEL ;
input [2:0] RXOUTCLKSEL ;
input [2:0] RXPRBSSEL ;
input [2:0] RXRATE ;
input [2:0] TXBUFDIFFCTRL ;
input [2:0] TXHEADER ;
input [2:0] TXMARGIN ;
input [2:0] TXOUTCLKSEL ;
input [2:0] TXPRBSSEL ;
input [2:0] TXRATE ;
input [31:0] TXDATA ;
input [3:0] RXCHBONDI ;
input [3:0] RXOSINTCFG ;
input [3:0] RXOSINTID0 ;
input [3:0] TX8B10BBYPASS ;
input [3:0] TXCHARDISPMODE ;
input [3:0] TXCHARDISPVAL ;
input [3:0] TXCHARISK ;
input [3:0] TXDIFFCTRL ;
input [4:0] TXPIPPMSTEPSIZE ;
input [4:0] TXPOSTCURSOR ;
input [4:0] TXPRECURSOR ;
input [6:0] TXMAINCURSOR ;
input [6:0] TXSEQUENCE ;
input [8:0] DRPADDR ;
output DRPRDY ;
output EYESCANDATAERROR ;
output GTPTXN ;
output GTPTXP ;
output PHYSTATUS ;
output PMARSVDOUT0 ;
output PMARSVDOUT1 ;
output RXBYTEISALIGNED ;
output RXBYTEREALIGN ;
output RXCDRLOCK ;
output RXCHANBONDSEQ ;
output RXCHANISALIGNED ;
output RXCHANREALIGN ;
output RXCOMINITDET ;
output RXCOMMADET ;
output RXCOMSASDET ;
output RXCOMWAKEDET ;
output RXDLYSRESETDONE ;
output RXELECIDLE ;
output RXHEADERVALID ;
output RXOSINTDONE ;
output RXOSINTSTARTED ;
output RXOSINTSTROBEDONE ;
output RXOSINTSTROBESTARTED ;
output RXOUTCLK ;
output RXOUTCLKFABRIC ;
output RXOUTCLKPCS ;
output RXPHALIGNDONE ;
output RXPMARESETDONE ;
output RXPRBSERR ;
output RXRATEDONE ;
output RXRESETDONE ;
output RXSYNCDONE ;
output RXSYNCOUT ;
output RXVALID ;
output TXCOMFINISH ;
output TXDLYSRESETDONE ;
output TXGEARBOXREADY ;
output TXOUTCLK ;
output TXOUTCLKFABRIC ;
output TXOUTCLKPCS ;
output TXPHALIGNDONE ;
output TXPHINITDONE ;
output TXPMARESETDONE ;
output TXRATEDONE ;
output TXRESETDONE ;
output TXSYNCDONE ;
output TXSYNCOUT ;
output [14:0] DMONITOROUT ;
output [15:0] DRPDO ;
output [15:0] PCSRSVDOUT ;
output [1:0] RXCLKCORCNT ;
output [1:0] RXDATAVALID ;
output [1:0] RXSTARTOFSEQ ;
output [1:0] TXBUFSTATUS ;
output [2:0] RXBUFSTATUS ;
output [2:0] RXHEADER ;
output [2:0] RXSTATUS ;
output [31:0] RXDATA ;
output [3:0] RXCHARISCOMMA ;
output [3:0] RXCHARISK ;
output [3:0] RXCHBONDO ;
output [3:0] RXDISPERR ;
output [3:0] RXNOTINTABLE ;
output [4:0] RXPHMONITOR ;
output [4:0] RXPHSLIPMONITOR ;
parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
parameter [0:0] ACJTAG_MODE = 1'b0;
parameter [0:0] ACJTAG_RESET = 1'b0;
parameter [19:0] ADAPT_CFG0 = 20'b00000000000000000000;
parameter ALIGN_COMMA_DOUBLE = "FALSE";
parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
parameter ALIGN_COMMA_WORD = 1;
parameter ALIGN_MCOMMA_DET = "TRUE";
parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
parameter ALIGN_PCOMMA_DET = "TRUE";
parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
parameter CBCC_DATA_SOURCE_SEL = "DECODED";
parameter [42:0] CFOK_CFG = 43'b1001001000000000000000001000000111010000000;
parameter [6:0] CFOK_CFG2 = 7'b0100000;
parameter [6:0] CFOK_CFG3 = 7'b0100000;
parameter [0:0] CFOK_CFG4 = 1'b0;
parameter [1:0] CFOK_CFG5 = 2'b00;
parameter [3:0] CFOK_CFG6 = 4'b0000;
parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
parameter CHAN_BOND_MAX_SKEW = 7;
parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
parameter CHAN_BOND_SEQ_2_USE = "FALSE";
parameter CHAN_BOND_SEQ_LEN = 1;
parameter [0:0] CLK_COMMON_SWING = 1'b0;
parameter CLK_CORRECT_USE = "TRUE";
parameter CLK_COR_KEEP_IDLE = "FALSE";
parameter CLK_COR_MAX_LAT = 20;
parameter CLK_COR_MIN_LAT = 18;
parameter CLK_COR_PRECEDENCE = "TRUE";
parameter CLK_COR_REPEAT_WAIT = 0;
parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
parameter CLK_COR_SEQ_2_USE = "FALSE";
parameter CLK_COR_SEQ_LEN = 1;
parameter DEC_MCOMMA_DETECT = "TRUE";
parameter DEC_PCOMMA_DETECT = "TRUE";
parameter DEC_VALID_COMMA_ONLY = "TRUE";
parameter [23:0] DMONITOR_CFG = 24'h000A00;
parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
parameter [5:0] ES_CONTROL = 6'b000000;
parameter ES_ERRDET_EN = "FALSE";
parameter ES_EYE_SCAN_EN = "FALSE";
parameter [11:0] ES_HORZ_OFFSET = 12'h010;
parameter [9:0] ES_PMA_CFG = 10'b0000000000;
parameter [4:0] ES_PRESCALE = 5'b00000;
parameter [79:0] ES_QUALIFIER = 80'h00000000000000000000;
parameter [79:0] ES_QUAL_MASK = 80'h00000000000000000000;
parameter [79:0] ES_SDATA_MASK = 80'h00000000000000000000;
parameter [8:0] ES_VERT_OFFSET = 9'b000000000;
parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
parameter FTS_LANE_DESKEW_EN = "FALSE";
parameter [2:0] GEARBOX_MODE = 3'b000;
parameter [0:0] LOOPBACK_CFG = 1'b0;
parameter [1:0] OUTREFCLK_SEL_INV = 2'b11;
parameter PCS_PCIE_EN = "FALSE";
parameter [47:0] PCS_RSVD_ATTR = 48'h000000000000;
parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
parameter [0:0] PMA_LOOPBACK_CFG = 1'b0;
parameter [31:0] PMA_RSV = 32'h00000333;
parameter [31:0] PMA_RSV2 = 32'h00002050;
parameter [1:0] PMA_RSV3 = 2'b00;
parameter [3:0] PMA_RSV4 = 4'b0000;
parameter [0:0] PMA_RSV5 = 1'b0;
parameter [0:0] PMA_RSV6 = 1'b0;
parameter [0:0] PMA_RSV7 = 1'b0;
parameter [4:0] RXBUFRESET_TIME = 5'b00001;
parameter RXBUF_ADDR_MODE = "FULL";
parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
parameter RXBUF_EN = "TRUE";
parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
parameter RXBUF_RESET_ON_EIDLE = "FALSE";
parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
parameter RXBUF_THRESH_OVFLW = 61;
parameter RXBUF_THRESH_OVRD = "FALSE";
parameter RXBUF_THRESH_UNDFLW = 4;
parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
parameter [82:0] RXCDR_CFG = 83'h0000107FE406001041010;
parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
parameter [5:0] RXCDR_LOCK_CFG = 6'b001001;
parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
parameter [15:0] RXDLY_CFG = 16'h0010;
parameter [8:0] RXDLY_LCFG = 9'h020;
parameter [15:0] RXDLY_TAP_CFG = 16'h0000;
parameter RXGEARBOX_EN = "FALSE";
parameter [4:0] RXISCANRESET_TIME = 5'b00001;
parameter [6:0] RXLPMRESET_TIME = 7'b0001111;
parameter [0:0] RXLPM_BIAS_STARTUP_DISABLE = 1'b0;
parameter [3:0] RXLPM_CFG = 4'b0110;
parameter [0:0] RXLPM_CFG1 = 1'b0;
parameter [0:0] RXLPM_CM_CFG = 1'b0;
parameter [8:0] RXLPM_GC_CFG = 9'b111100010;
parameter [2:0] RXLPM_GC_CFG2 = 3'b001;
parameter [13:0] RXLPM_HF_CFG = 14'b00001111110000;
parameter [4:0] RXLPM_HF_CFG2 = 5'b01010;
parameter [3:0] RXLPM_HF_CFG3 = 4'b0000;
parameter [0:0] RXLPM_HOLD_DURING_EIDLE = 1'b0;
parameter [0:0] RXLPM_INCM_CFG = 1'b0;
parameter [0:0] RXLPM_IPCM_CFG = 1'b0;
parameter [17:0] RXLPM_LF_CFG = 18'b000000001111110000;
parameter [4:0] RXLPM_LF_CFG2 = 5'b01010;
parameter [2:0] RXLPM_OSINT_CFG = 3'b100;
parameter [6:0] RXOOB_CFG = 7'b0000110;
parameter RXOOB_CLK_CFG = "PMA";
parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
parameter [4:0] RXOSCALRESET_TIMEOUT = 5'b00000;
parameter RXOUT_DIV = 2;
parameter [4:0] RXPCSRESET_TIME = 5'b00001;
parameter [23:0] RXPHDLY_CFG = 24'h084000;
parameter [23:0] RXPH_CFG = 24'hC00002;
parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
parameter [2:0] RXPI_CFG0 = 3'b000;
parameter [0:0] RXPI_CFG1 = 1'b0;
parameter [0:0] RXPI_CFG2 = 1'b0;
parameter [4:0] RXPMARESET_TIME = 5'b00011;
parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
parameter RXSLIDE_AUTO_WAIT = 7;
parameter RXSLIDE_MODE = "OFF";
parameter [0:0] RXSYNC_MULTILANE = 1'b0;
parameter [0:0] RXSYNC_OVRD = 1'b0;
parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
parameter [15:0] RX_BIAS_CFG = 16'b0000111100110011;
parameter [5:0] RX_BUFFER_CFG = 6'b000000;
parameter RX_CLK25_DIV = 7;
parameter [0:0] RX_CLKMUX_EN = 1'b1;
parameter [1:0] RX_CM_SEL = 2'b11;
parameter [3:0] RX_CM_TRIM = 4'b0100;
parameter RX_DATA_WIDTH = 20;
parameter [5:0] RX_DDI_SEL = 6'b000000;
parameter [13:0] RX_DEBUG_CFG = 14'b00000000000000;
parameter RX_DEFER_RESET_BUF_EN = "TRUE";
parameter RX_DISPERR_SEQ_MATCH = "TRUE";
parameter [12:0] RX_OS_CFG = 13'b0001111110000;
parameter RX_SIG_VALID_DLY = 10;
parameter RX_XCLK_SEL = "RXREC";
parameter SAS_MAX_COM = 64;
parameter SAS_MIN_COM = 36;
parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
parameter [2:0] SATA_BURST_VAL = 3'b100;
parameter [2:0] SATA_EIDLE_VAL = 3'b100;
parameter SATA_MAX_BURST = 8;
parameter SATA_MAX_INIT = 21;
parameter SATA_MAX_WAKE = 7;
parameter SATA_MIN_BURST = 4;
parameter SATA_MIN_INIT = 12;
parameter SATA_MIN_WAKE = 4;
parameter SATA_PLL_CFG = "VCO_3000MHZ";
parameter SHOW_REALIGN_COMMA = "TRUE";
parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
parameter SIM_RESET_SPEEDUP = "TRUE";
parameter SIM_TX_EIDLE_DRIVE_LEVEL = "X";
parameter SIM_VERSION = "1.0";
parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
parameter [2:0] TERM_RCAL_OVRD = 3'b000;
parameter [7:0] TRANS_TIME_RATE = 8'h0E;
parameter [31:0] TST_RSV = 32'h00000000;
parameter TXBUF_EN = "TRUE";
parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
parameter [15:0] TXDLY_CFG = 16'h0010;
parameter [8:0] TXDLY_LCFG = 9'h020;
parameter [15:0] TXDLY_TAP_CFG = 16'h0000;
parameter TXGEARBOX_EN = "FALSE";
parameter [0:0] TXOOB_CFG = 1'b0;
parameter TXOUT_DIV = 2;
parameter [4:0] TXPCSRESET_TIME = 5'b00001;
parameter [23:0] TXPHDLY_CFG = 24'h084000;
parameter [15:0] TXPH_CFG = 16'h0400;
parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
parameter [1:0] TXPI_CFG0 = 2'b00;
parameter [1:0] TXPI_CFG1 = 2'b00;
parameter [1:0] TXPI_CFG2 = 2'b00;
parameter [0:0] TXPI_CFG3 = 1'b0;
parameter [0:0] TXPI_CFG4 = 1'b0;
parameter [2:0] TXPI_CFG5 = 3'b000;
parameter [0:0] TXPI_GREY_SEL = 1'b0;
parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
parameter TXPI_PPMCLK_SEL = "TXUSRCLK2";
parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
parameter [4:0] TXPMARESET_TIME = 5'b00001;
parameter [0:0] TXSYNC_MULTILANE = 1'b0;
parameter [0:0] TXSYNC_OVRD = 1'b0;
parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
parameter TX_CLK25_DIV = 7;
parameter [0:0] TX_CLKMUX_EN = 1'b1;
parameter TX_DATA_WIDTH = 20;
parameter [5:0] TX_DEEMPH0 = 6'b000000;
parameter [5:0] TX_DEEMPH1 = 6'b000000;
parameter TX_DRIVE_MODE = "DIRECT";
parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
parameter [0:0] TX_PREDRIVER_MODE = 1'b0;
parameter [13:0] TX_RXDETECT_CFG = 14'h1832;
parameter [2:0] TX_RXDETECT_REF = 3'b100;
parameter TX_XCLK_SEL = "TXUSR";
parameter [0:0] UCODEER_CLR = 1'b0;
parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: GTPE2_CHANNEL ####

//#### BEGIN MODULE DEFINITION FOR :GTPE2_COMMON ###
module GTPE2_COMMON (
  DMONITOROUT,
  DRPDO,
  DRPRDY,
  PLL0FBCLKLOST,
  PLL0LOCK,
  PLL0OUTCLK,
  PLL0OUTREFCLK,
  PLL0REFCLKLOST,
  PLL1FBCLKLOST,
  PLL1LOCK,
  PLL1OUTCLK,
  PLL1OUTREFCLK,
  PLL1REFCLKLOST,
  PMARSVDOUT,
  REFCLKOUTMONITOR0,
  REFCLKOUTMONITOR1,

  BGBYPASSB,
  BGMONITORENB,
  BGPDB,
  BGRCALOVRD,
  BGRCALOVRDENB,
  DRPADDR,
  DRPCLK,
  DRPDI,
  DRPEN,
  DRPWE,
  GTEASTREFCLK0,
  GTEASTREFCLK1,
  GTGREFCLK0,
  GTGREFCLK1,
  GTREFCLK0,
  GTREFCLK1,
  GTWESTREFCLK0,
  GTWESTREFCLK1,
  PLL0LOCKDETCLK,
  PLL0LOCKEN,
  PLL0PD,
  PLL0REFCLKSEL,
  PLL0RESET,
  PLL1LOCKDETCLK,
  PLL1LOCKEN,
  PLL1PD,
  PLL1REFCLKSEL,
  PLL1RESET,
  PLLRSVD1,
  PLLRSVD2,
  PMARSVD,
  RCALENB
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input BGBYPASSB ;
input BGMONITORENB ;
input BGPDB ;
input BGRCALOVRDENB ;
input DRPCLK ;
input DRPEN ;
input DRPWE ;
input GTEASTREFCLK0 ;
input GTEASTREFCLK1 ;
input GTGREFCLK0 ;
input GTGREFCLK1 ;
input GTREFCLK0 ;
input GTREFCLK1 ;
input GTWESTREFCLK0 ;
input GTWESTREFCLK1 ;
input PLL0LOCKDETCLK ;
input PLL0LOCKEN ;
input PLL0PD ;
input PLL0RESET ;
input PLL1LOCKDETCLK ;
input PLL1LOCKEN ;
input PLL1PD ;
input PLL1RESET ;
input RCALENB ;
input [15:0] DRPDI ;
input [15:0] PLLRSVD1 ;
input [2:0] PLL0REFCLKSEL ;
input [2:0] PLL1REFCLKSEL ;
input [4:0] BGRCALOVRD ;
input [4:0] PLLRSVD2 ;
input [7:0] DRPADDR ;
input [7:0] PMARSVD ;
output DRPRDY ;
output PLL0FBCLKLOST ;
output PLL0LOCK ;
output PLL0OUTCLK ;
output PLL0OUTREFCLK ;
output PLL0REFCLKLOST ;
output PLL1FBCLKLOST ;
output PLL1LOCK ;
output PLL1OUTCLK ;
output PLL1OUTREFCLK ;
output PLL1REFCLKLOST ;
output REFCLKOUTMONITOR0 ;
output REFCLKOUTMONITOR1 ;
output [15:0] DRPDO ;
output [15:0] PMARSVDOUT ;
output [7:0] DMONITOROUT ;
parameter [63:0] BIAS_CFG = 64'h0000000000000000;
parameter [31:0] COMMON_CFG = 32'h00000000;
parameter [26:0] PLL0_CFG = 27'h01F03DC;
parameter [0:0] PLL0_DMON_CFG = 1'b0;
parameter PLL0_FBDIV = 4;
parameter PLL0_FBDIV_45 = 5;
parameter [23:0] PLL0_INIT_CFG = 24'h00001E;
parameter [8:0] PLL0_LOCK_CFG = 9'h1E8;
parameter PLL0_REFCLK_DIV = 1;
parameter [26:0] PLL1_CFG = 27'h01F03DC;
parameter [0:0] PLL1_DMON_CFG = 1'b0;
parameter PLL1_FBDIV = 4;
parameter PLL1_FBDIV_45 = 5;
parameter [23:0] PLL1_INIT_CFG = 24'h00001E;
parameter [8:0] PLL1_LOCK_CFG = 9'h1E8;
parameter PLL1_REFCLK_DIV = 1;
parameter [7:0] PLL_CLKOUT_CFG = 8'b00000000;
parameter [15:0] RSVD_ATTR0 = 16'h0000;
parameter [15:0] RSVD_ATTR1 = 16'h0000;
parameter [2:0] SIM_PLL0REFCLK_SEL = 3'b001;
parameter [2:0] SIM_PLL1REFCLK_SEL = 3'b001;
parameter SIM_RESET_SPEEDUP = "TRUE";
parameter SIM_VERSION = "1.0";
endmodule
//#### END MODULE DEFINITION FOR: GTPE2_COMMON ####

//#### BEGIN MODULE DEFINITION FOR :GTP_DUAL ###
module GTP_DUAL (
	DO,
	DRDY,
	PHYSTATUS0,
	PHYSTATUS1,
	PLLLKDET,
	REFCLKOUT,
	RESETDONE0,
	RESETDONE1,
	RXBUFSTATUS0,
	RXBUFSTATUS1,
	RXBYTEISALIGNED0,
	RXBYTEISALIGNED1,
	RXBYTEREALIGN0,
	RXBYTEREALIGN1,
	RXCHANBONDSEQ0,
	RXCHANBONDSEQ1,
	RXCHANISALIGNED0,
	RXCHANISALIGNED1,
	RXCHANREALIGN0,
	RXCHANREALIGN1,
	RXCHARISCOMMA0,
	RXCHARISCOMMA1,
	RXCHARISK0,
	RXCHARISK1,
	RXCHBONDO0,
	RXCHBONDO1,
	RXCLKCORCNT0,
	RXCLKCORCNT1,
	RXCOMMADET0,
	RXCOMMADET1,
	RXDATA0,
	RXDATA1,
	RXDISPERR0,
	RXDISPERR1,
	RXELECIDLE0,
	RXELECIDLE1,
	RXLOSSOFSYNC0,
	RXLOSSOFSYNC1,
	RXNOTINTABLE0,
	RXNOTINTABLE1,
	RXOVERSAMPLEERR0,
	RXOVERSAMPLEERR1,
	RXPRBSERR0,
	RXPRBSERR1,
	RXRECCLK0,
	RXRECCLK1,
	RXRUNDISP0,
	RXRUNDISP1,
	RXSTATUS0,
	RXSTATUS1,
	RXVALID0,
	RXVALID1,
	TXBUFSTATUS0,
	TXBUFSTATUS1,
	TXKERR0,
	TXKERR1,
	TXN0,
	TXN1,
	TXOUTCLK0,
	TXOUTCLK1,
	TXP0,
	TXP1,
	TXRUNDISP0,
	TXRUNDISP1,

	CLKIN,
	DADDR,
	DCLK,
	DEN,
	DI,
	DWE,
	GTPRESET,
	GTPTEST,
	INTDATAWIDTH,
	LOOPBACK0,
	LOOPBACK1,
	PLLLKDETEN,
	PLLPOWERDOWN,
	PRBSCNTRESET0,
	PRBSCNTRESET1,
	REFCLKPWRDNB,
	RXBUFRESET0,
	RXBUFRESET1,
	RXCDRRESET0,
	RXCDRRESET1,
	RXCHBONDI0,
	RXCHBONDI1,
	RXCOMMADETUSE0,
	RXCOMMADETUSE1,
	RXDATAWIDTH0,
	RXDATAWIDTH1,
	RXDEC8B10BUSE0,
	RXDEC8B10BUSE1,
	RXELECIDLERESET0,
	RXELECIDLERESET1,	 
	RXENCHANSYNC0,
	RXENCHANSYNC1,
        RXENELECIDLERESETB,	 
	RXENEQB0,
	RXENEQB1,
	RXENMCOMMAALIGN0,
	RXENMCOMMAALIGN1,
	RXENPCOMMAALIGN0,
	RXENPCOMMAALIGN1,
	RXENPRBSTST0,
	RXENPRBSTST1,
	RXENSAMPLEALIGN0,
	RXENSAMPLEALIGN1,
	RXEQMIX0,
	RXEQMIX1,
	RXEQPOLE0,
	RXEQPOLE1,
	RXN0,
	RXN1,
	RXP0,
	RXP1,
	RXPMASETPHASE0,
	RXPMASETPHASE1,
	RXPOLARITY0,
	RXPOLARITY1,
	RXPOWERDOWN0,
	RXPOWERDOWN1,
	RXRESET0,
	RXRESET1,
	RXSLIDE0,
	RXSLIDE1,
	RXUSRCLK0,
	RXUSRCLK1,
	RXUSRCLK20,
	RXUSRCLK21,
	TXBUFDIFFCTRL0,
	TXBUFDIFFCTRL1,
	TXBYPASS8B10B0,
	TXBYPASS8B10B1,
	TXCHARDISPMODE0,
	TXCHARDISPMODE1,
	TXCHARDISPVAL0,
	TXCHARDISPVAL1,
	TXCHARISK0,
	TXCHARISK1,
	TXCOMSTART0,
	TXCOMSTART1,
	TXCOMTYPE0,
	TXCOMTYPE1,
	TXDATA0,
	TXDATA1,
	TXDATAWIDTH0,
	TXDATAWIDTH1,
	TXDETECTRX0,
	TXDETECTRX1,
	TXDIFFCTRL0,
	TXDIFFCTRL1,
	TXELECIDLE0,
	TXELECIDLE1,
	TXENC8B10BUSE0,
	TXENC8B10BUSE1,
	TXENPMAPHASEALIGN,
	TXENPRBSTST0,
	TXENPRBSTST1,
	TXINHIBIT0,
	TXINHIBIT1,
	TXPMASETPHASE,
	TXPOLARITY0,
	TXPOLARITY1,
	TXPOWERDOWN0,
	TXPOWERDOWN1,
	TXPREEMPHASIS0,
	TXPREEMPHASIS1,
	TXRESET0,
	TXRESET1,
	TXUSRCLK0,
	TXUSRCLK1,
	TXUSRCLK20,
	TXUSRCLK21

) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKIN ;
input DCLK ;
input DEN ;
input DWE ;
input GTPRESET ;
input INTDATAWIDTH ;
input PLLLKDETEN ;
input PLLPOWERDOWN ;
input PRBSCNTRESET0 ;
input PRBSCNTRESET1 ;
input REFCLKPWRDNB ;
input RXBUFRESET0 ;
input RXBUFRESET1 ;
input RXCDRRESET0 ;
input RXCDRRESET1 ;
input RXCOMMADETUSE0 ;
input RXCOMMADETUSE1 ;
input RXDATAWIDTH0 ;
input RXDATAWIDTH1 ;
input RXDEC8B10BUSE0 ;
input RXDEC8B10BUSE1 ;
input RXELECIDLERESET0 ;
input RXELECIDLERESET1 ;
input RXENCHANSYNC0 ;
input RXENCHANSYNC1 ;
input RXENELECIDLERESETB ;
input RXENEQB0 ;
input RXENEQB1 ;
input RXENMCOMMAALIGN0 ;
input RXENMCOMMAALIGN1 ;
input RXENPCOMMAALIGN0 ;
input RXENPCOMMAALIGN1 ;
input RXENSAMPLEALIGN0 ;
input RXENSAMPLEALIGN1 ;
input RXN0 ;
input RXN1 ;
input RXP0 ;
input RXP1 ;
input RXPMASETPHASE0 ;
input RXPMASETPHASE1 ;
input RXPOLARITY0 ;
input RXPOLARITY1 ;
input RXRESET0 ;
input RXRESET1 ;
input RXSLIDE0 ;
input RXSLIDE1 ;
input RXUSRCLK0 ;
input RXUSRCLK1 ;
input RXUSRCLK20 ;
input RXUSRCLK21 ;
input TXCOMSTART0 ;
input TXCOMSTART1 ;
input TXCOMTYPE0 ;
input TXCOMTYPE1 ;
input TXDATAWIDTH0 ;
input TXDATAWIDTH1 ;
input TXDETECTRX0 ;
input TXDETECTRX1 ;
input TXELECIDLE0 ;
input TXELECIDLE1 ;
input TXENC8B10BUSE0 ;
input TXENC8B10BUSE1 ;
input TXENPMAPHASEALIGN ;
input TXINHIBIT0 ;
input TXINHIBIT1 ;
input TXPMASETPHASE ;
input TXPOLARITY0 ;
input TXPOLARITY1 ;
input TXRESET0 ;
input TXRESET1 ;
input TXUSRCLK0 ;
input TXUSRCLK1 ;
input TXUSRCLK20 ;
input TXUSRCLK21 ;
input [15:0] DI ;
input [15:0] TXDATA0 ;
input [15:0] TXDATA1 ;
input [1:0] RXENPRBSTST0 ;
input [1:0] RXENPRBSTST1 ;
input [1:0] RXEQMIX0 ;
input [1:0] RXEQMIX1 ;
input [1:0] RXPOWERDOWN0 ;
input [1:0] RXPOWERDOWN1 ;
input [1:0] TXBYPASS8B10B0 ;
input [1:0] TXBYPASS8B10B1 ;
input [1:0] TXCHARDISPMODE0 ;
input [1:0] TXCHARDISPMODE1 ;
input [1:0] TXCHARDISPVAL0 ;
input [1:0] TXCHARDISPVAL1 ;
input [1:0] TXCHARISK0 ;
input [1:0] TXCHARISK1 ;
input [1:0] TXENPRBSTST0 ;
input [1:0] TXENPRBSTST1 ;
input [1:0] TXPOWERDOWN0 ;
input [1:0] TXPOWERDOWN1 ;
input [2:0] LOOPBACK0 ;
input [2:0] LOOPBACK1 ;
input [2:0] RXCHBONDI0 ;
input [2:0] RXCHBONDI1 ;
input [2:0] TXBUFDIFFCTRL0 ;
input [2:0] TXBUFDIFFCTRL1 ;
input [2:0] TXDIFFCTRL0 ;
input [2:0] TXDIFFCTRL1 ;
input [2:0] TXPREEMPHASIS0 ;
input [2:0] TXPREEMPHASIS1 ;
input [3:0] GTPTEST ;
input [3:0] RXEQPOLE0 ;
input [3:0] RXEQPOLE1 ;
input [6:0] DADDR ;
output DRDY ;
output PHYSTATUS0 ;
output PHYSTATUS1 ;
output PLLLKDET ;
output REFCLKOUT ;
output RESETDONE0 ;
output RESETDONE1 ;
output RXBYTEISALIGNED0 ;
output RXBYTEISALIGNED1 ;
output RXBYTEREALIGN0 ;
output RXBYTEREALIGN1 ;
output RXCHANBONDSEQ0 ;
output RXCHANBONDSEQ1 ;
output RXCHANISALIGNED0 ;
output RXCHANISALIGNED1 ;
output RXCHANREALIGN0 ;
output RXCHANREALIGN1 ;
output RXCOMMADET0 ;
output RXCOMMADET1 ;
output RXELECIDLE0 ;
output RXELECIDLE1 ;
output RXOVERSAMPLEERR0 ;
output RXOVERSAMPLEERR1 ;
output RXPRBSERR0 ;
output RXPRBSERR1 ;
output RXRECCLK0 ;
output RXRECCLK1 ;
output RXVALID0 ;
output RXVALID1 ;
output TXN0 ;
output TXN1 ;
output TXOUTCLK0 ;
output TXOUTCLK1 ;
output TXP0 ;
output TXP1 ;
output [15:0] DO ;
output [15:0] RXDATA0 ;
output [15:0] RXDATA1 ;
output [1:0] RXCHARISCOMMA0 ;
output [1:0] RXCHARISCOMMA1 ;
output [1:0] RXCHARISK0 ;
output [1:0] RXCHARISK1 ;
output [1:0] RXDISPERR0 ;
output [1:0] RXDISPERR1 ;
output [1:0] RXLOSSOFSYNC0 ;
output [1:0] RXLOSSOFSYNC1 ;
output [1:0] RXNOTINTABLE0 ;
output [1:0] RXNOTINTABLE1 ;
output [1:0] RXRUNDISP0 ;
output [1:0] RXRUNDISP1 ;
output [1:0] TXBUFSTATUS0 ;
output [1:0] TXBUFSTATUS1 ;
output [1:0] TXKERR0 ;
output [1:0] TXKERR1 ;
output [1:0] TXRUNDISP0 ;
output [1:0] TXRUNDISP1 ;
output [2:0] RXBUFSTATUS0 ;
output [2:0] RXBUFSTATUS1 ;
output [2:0] RXCHBONDO0 ;
output [2:0] RXCHBONDO1 ;
output [2:0] RXCLKCORCNT0 ;
output [2:0] RXCLKCORCNT1 ;
output [2:0] RXSTATUS0 ;
output [2:0] RXSTATUS1 ;
parameter AC_CAP_DIS_0 = "TRUE";
parameter AC_CAP_DIS_1 = "TRUE";
parameter CHAN_BOND_MODE_0 = "OFF";
parameter CHAN_BOND_MODE_1 = "OFF";
parameter CHAN_BOND_SEQ_2_USE_0 = "TRUE";
parameter CHAN_BOND_SEQ_2_USE_1 = "TRUE";
parameter CLKINDC_B = "TRUE";
parameter CLK_CORRECT_USE_0 = "TRUE";
parameter CLK_CORRECT_USE_1 = "TRUE";
parameter CLK_COR_INSERT_IDLE_FLAG_0 = "FALSE";
parameter CLK_COR_INSERT_IDLE_FLAG_1 = "FALSE";
parameter CLK_COR_KEEP_IDLE_0 = "FALSE";
parameter CLK_COR_KEEP_IDLE_1 = "FALSE";
parameter CLK_COR_PRECEDENCE_0 = "TRUE";
parameter CLK_COR_PRECEDENCE_1 = "TRUE";
parameter CLK_COR_SEQ_2_USE_0 = "FALSE";
parameter CLK_COR_SEQ_2_USE_1 = "FALSE";
parameter COMMA_DOUBLE_0 = "FALSE";
parameter COMMA_DOUBLE_1 = "FALSE";
parameter DEC_MCOMMA_DETECT_0 = "TRUE";
parameter DEC_MCOMMA_DETECT_1 = "TRUE";
parameter DEC_PCOMMA_DETECT_0 = "TRUE";
parameter DEC_PCOMMA_DETECT_1 = "TRUE";
parameter DEC_VALID_COMMA_ONLY_0 = "TRUE";
parameter DEC_VALID_COMMA_ONLY_1 = "TRUE";
parameter MCOMMA_DETECT_0 = "TRUE";
parameter MCOMMA_DETECT_1 = "TRUE";
parameter OVERSAMPLE_MODE = "FALSE";
parameter PCI_EXPRESS_MODE_0 = "TRUE";
parameter PCI_EXPRESS_MODE_1 = "TRUE";
parameter PCOMMA_DETECT_0 = "TRUE";
parameter PCOMMA_DETECT_1 = "TRUE";
parameter PLL_SATA_0 = "FALSE";
parameter PLL_SATA_1 = "FALSE";
parameter RCV_TERM_GND_0 = "TRUE";
parameter RCV_TERM_GND_1 = "TRUE";
parameter RCV_TERM_MID_0 = "FALSE";
parameter RCV_TERM_MID_1 = "FALSE";
parameter RCV_TERM_VTTRX_0 = "FALSE";
parameter RCV_TERM_VTTRX_1 = "FALSE";
parameter RX_BUFFER_USE_0 = "TRUE";
parameter RX_BUFFER_USE_1 = "TRUE";
parameter RX_DECODE_SEQ_MATCH_0 = "TRUE";
parameter RX_DECODE_SEQ_MATCH_1 = "TRUE";
parameter RX_LOSS_OF_SYNC_FSM_0 = "FALSE";
parameter RX_LOSS_OF_SYNC_FSM_1 = "FALSE";
parameter RX_SLIDE_MODE_0 = "PCS";
parameter RX_SLIDE_MODE_1 = "PCS";
parameter RX_STATUS_FMT_0 = "PCIE";
parameter RX_STATUS_FMT_1 = "PCIE";
parameter RX_XCLK_SEL_0 = "RXREC";
parameter RX_XCLK_SEL_1 = "RXREC";
parameter SIM_MODE = "FAST";
parameter SIM_PLL_PERDIV2 = 9'h190;
parameter SIM_RECEIVER_DETECT_PASS0 = "FALSE";
parameter SIM_RECEIVER_DETECT_PASS1 = "FALSE";
parameter TERMINATION_OVRD = "FALSE";
parameter TX_BUFFER_USE_0 = "TRUE";
parameter TX_BUFFER_USE_1 = "TRUE";
parameter TX_DIFF_BOOST_0 = "TRUE";
parameter TX_DIFF_BOOST_1 = "TRUE";
parameter TX_XCLK_SEL_0 = "TXUSR";
parameter TX_XCLK_SEL_1 = "TXUSR";
parameter [15:0] TRANS_TIME_FROM_P2_0 = 16'h003c;
parameter [15:0] TRANS_TIME_FROM_P2_1 = 16'h003c;
parameter [15:0] TRANS_TIME_NON_P2_0 = 16'h0019;
parameter [15:0] TRANS_TIME_NON_P2_1 = 16'h0019;
parameter [15:0] TRANS_TIME_TO_P2_0 = 16'h0064;
parameter [15:0] TRANS_TIME_TO_P2_1 = 16'h0064;
parameter [24:0] PMA_RX_CFG_0 = 25'h09f0089;
parameter [24:0] PMA_RX_CFG_1 = 25'h09f0089;
parameter [26:0] PMA_CDR_SCAN_0 = 27'h6c07640;
parameter [26:0] PMA_CDR_SCAN_1 = 27'h6c07640;
parameter [27:0] PCS_COM_CFG = 28'h1680a0e;
parameter [2:0] OOBDETECT_THRESHOLD_0 = 3'b001;
parameter [2:0] OOBDETECT_THRESHOLD_1 = 3'b001;
parameter [2:0] SATA_BURST_VAL_0 = 3'b100;
parameter [2:0] SATA_BURST_VAL_1 = 3'b100;
parameter [2:0] SATA_IDLE_VAL_0 = 3'b011;
parameter [2:0] SATA_IDLE_VAL_1 = 3'b011;
parameter [31:0] PRBS_ERR_THRESHOLD_0 = 32'h1;
parameter [31:0] PRBS_ERR_THRESHOLD_1 = 32'h1;
parameter [3:0] CHAN_BOND_SEQ_1_ENABLE_0 = 4'b1111;
parameter [3:0] CHAN_BOND_SEQ_1_ENABLE_1 = 4'b1111;
parameter [3:0] CHAN_BOND_SEQ_2_ENABLE_0 = 4'b1111;
parameter [3:0] CHAN_BOND_SEQ_2_ENABLE_1 = 4'b1111;
parameter [3:0] CLK_COR_SEQ_1_ENABLE_0 = 4'b1111;
parameter [3:0] CLK_COR_SEQ_1_ENABLE_1 = 4'b1111;
parameter [3:0] CLK_COR_SEQ_2_ENABLE_0 = 4'b1111;
parameter [3:0] CLK_COR_SEQ_2_ENABLE_1 = 4'b1111;
parameter [3:0] COM_BURST_VAL_0 = 4'b1111;
parameter [3:0] COM_BURST_VAL_1 = 4'b1111;
parameter [4:0] TERMINATION_CTRL = 5'b10100;
parameter [4:0] TXRX_INVERT_0 = 5'b00000;
parameter [4:0] TXRX_INVERT_1 = 5'b00000;
parameter [9:0] CHAN_BOND_SEQ_1_1_0 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_1_1 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_2_0 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_2_1 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_3_0 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_3_1 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_4_0 = 10'b0110111100;
parameter [9:0] CHAN_BOND_SEQ_1_4_1 = 10'b0110111100;
parameter [9:0] CHAN_BOND_SEQ_2_1_0 = 10'b0110111100;
parameter [9:0] CHAN_BOND_SEQ_2_1_1 = 10'b0110111100;
parameter [9:0] CHAN_BOND_SEQ_2_2_0 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_2_1 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_3_0 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_3_1 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_4_0 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_4_1 = 10'b0100111100;
parameter [9:0] CLK_COR_SEQ_1_1_0 = 10'b0100011100;
parameter [9:0] CLK_COR_SEQ_1_1_1 = 10'b0100011100;
parameter [9:0] CLK_COR_SEQ_1_2_0 = 10'b0;
parameter [9:0] CLK_COR_SEQ_1_2_1 = 10'b0;
parameter [9:0] CLK_COR_SEQ_1_3_0 = 10'b0;
parameter [9:0] CLK_COR_SEQ_1_3_1 = 10'b0;
parameter [9:0] CLK_COR_SEQ_1_4_0 = 10'b0;
parameter [9:0] CLK_COR_SEQ_1_4_1 = 10'b0;
parameter [9:0] CLK_COR_SEQ_2_1_0 = 10'b0;
parameter [9:0] CLK_COR_SEQ_2_1_1 = 10'b0;
parameter [9:0] CLK_COR_SEQ_2_2_0 = 10'b0;
parameter [9:0] CLK_COR_SEQ_2_2_1 = 10'b0;
parameter [9:0] CLK_COR_SEQ_2_3_0 = 10'b0;
parameter [9:0] CLK_COR_SEQ_2_3_1 = 10'b0;
parameter [9:0] CLK_COR_SEQ_2_4_0 = 10'b0;
parameter [9:0] CLK_COR_SEQ_2_4_1 = 10'b0;
parameter [9:0] COMMA_10B_ENABLE_0 = 10'b1111111111;
parameter [9:0] COMMA_10B_ENABLE_1 = 10'b1111111111;
parameter [9:0] MCOMMA_10B_VALUE_0 = 10'b1010000011;
parameter [9:0] MCOMMA_10B_VALUE_1 = 10'b1010000011;
parameter [9:0] PCOMMA_10B_VALUE_0 = 10'b0101111100;
parameter [9:0] PCOMMA_10B_VALUE_1 = 10'b0101111100;
parameter ALIGN_COMMA_WORD_0 = 1;
parameter ALIGN_COMMA_WORD_1 = 1;
parameter CHAN_BOND_1_MAX_SKEW_0 = 7;
parameter CHAN_BOND_1_MAX_SKEW_1 = 7;
parameter CHAN_BOND_2_MAX_SKEW_0 = 1;
parameter CHAN_BOND_2_MAX_SKEW_1 = 1;
parameter CHAN_BOND_LEVEL_0 = 0;
parameter CHAN_BOND_LEVEL_1 = 0;
parameter CHAN_BOND_SEQ_LEN_0 = 4;
parameter CHAN_BOND_SEQ_LEN_1 = 4;
parameter CLK25_DIVIDER = 4;
parameter CLK_COR_ADJ_LEN_0 = 1;
parameter CLK_COR_ADJ_LEN_1 = 1;
parameter CLK_COR_DET_LEN_0 = 1;
parameter CLK_COR_DET_LEN_1 = 1;
parameter CLK_COR_MAX_LAT_0 = 18;
parameter CLK_COR_MAX_LAT_1 = 18;
parameter CLK_COR_MIN_LAT_0 = 16;
parameter CLK_COR_MIN_LAT_1 = 16;
parameter CLK_COR_REPEAT_WAIT_0 = 5;
parameter CLK_COR_REPEAT_WAIT_1 = 5;
parameter OOB_CLK_DIVIDER = 4;
parameter PLL_DIVSEL_FB = 5;
parameter PLL_DIVSEL_REF = 2;
parameter PLL_RXDIVSEL_OUT_0 = 1;
parameter PLL_RXDIVSEL_OUT_1 = 1;
parameter PLL_TXDIVSEL_COMM_OUT = 1;
parameter PLL_TXDIVSEL_OUT_0 = 1;
parameter PLL_TXDIVSEL_OUT_1 = 1;
parameter RX_LOS_INVALID_INCR_0 = 8;
parameter RX_LOS_INVALID_INCR_1 = 8;
parameter RX_LOS_THRESHOLD_0 = 128;
parameter RX_LOS_THRESHOLD_1 = 128;
parameter SATA_MAX_BURST_0 = 7;
parameter SATA_MAX_BURST_1 = 7;
parameter SATA_MAX_INIT_0 = 22;
parameter SATA_MAX_INIT_1 = 22;
parameter SATA_MAX_WAKE_0 = 7;
parameter SATA_MAX_WAKE_1 = 7;
parameter SATA_MIN_BURST_0 = 4;
parameter SATA_MIN_BURST_1 = 4;
parameter SATA_MIN_INIT_0 = 12;
parameter SATA_MIN_INIT_1 = 12;
parameter SATA_MIN_WAKE_0 = 4;
parameter SATA_MIN_WAKE_1 = 4;
parameter SIM_GTPRESET_SPEEDUP = 0;
parameter TERMINATION_IMP_0 = 50;
parameter TERMINATION_IMP_1 = 50;
parameter TX_SYNC_FILTERB = 1;
endmodule
//#### END MODULE DEFINITION FOR: GTP_DUAL ####

//#### BEGIN MODULE DEFINITION FOR :GTXE1 ###
module GTXE1 (
  COMFINISH,
  COMINITDET,
  COMSASDET,
  COMWAKEDET,
  DFECLKDLYADJMON,
  DFEEYEDACMON,
  DFESENSCAL,
  DFETAP1MONITOR,
  DFETAP2MONITOR,
  DFETAP3MONITOR,
  DFETAP4MONITOR,
  DRDY,
  DRPDO,
  MGTREFCLKFAB,
  PHYSTATUS,
  RXBUFSTATUS,
  RXBYTEISALIGNED,
  RXBYTEREALIGN,
  RXCHANBONDSEQ,
  RXCHANISALIGNED,
  RXCHANREALIGN,
  RXCHARISCOMMA,
  RXCHARISK,
  RXCHBONDO,
  RXCLKCORCNT,
  RXCOMMADET,
  RXDATA,
  RXDATAVALID,
  RXDISPERR,
  RXDLYALIGNMONITOR,
  RXELECIDLE,
  RXHEADER,
  RXHEADERVALID,
  RXLOSSOFSYNC,
  RXNOTINTABLE,
  RXOVERSAMPLEERR,
  RXPLLLKDET,
  RXPRBSERR,
  RXRATEDONE,
  RXRECCLK,
  RXRECCLKPCS,
  RXRESETDONE,
  RXRUNDISP,
  RXSTARTOFSEQ,
  RXSTATUS,
  RXVALID,
  TSTOUT,
  TXBUFSTATUS,
  TXDLYALIGNMONITOR,
  TXGEARBOXREADY,
  TXKERR,
  TXN,
  TXOUTCLK,
  TXOUTCLKPCS,
  TXP,
  TXPLLLKDET,
  TXRATEDONE,
  TXRESETDONE,
  TXRUNDISP,
  DADDR,
  DCLK,
  DEN,
  DFECLKDLYADJ,
  DFEDLYOVRD,
  DFETAP1,
  DFETAP2,
  DFETAP3,
  DFETAP4,
  DFETAPOVRD,
  DI,
  DWE,
  GATERXELECIDLE,
  GREFCLKRX,
  GREFCLKTX,
  GTXRXRESET,
  GTXTEST,
  GTXTXRESET,
  IGNORESIGDET,
  LOOPBACK,
  MGTREFCLKRX,
  MGTREFCLKTX,
  NORTHREFCLKRX,
  NORTHREFCLKTX,
  PERFCLKRX,
  PERFCLKTX,
  PLLRXRESET,
  PLLTXRESET,
  PRBSCNTRESET,
  RXBUFRESET,
  RXCDRRESET,
  RXCHBONDI,
  RXCHBONDLEVEL,
  RXCHBONDMASTER,
  RXCHBONDSLAVE,
  RXCOMMADETUSE,
  RXDEC8B10BUSE,
  RXDLYALIGNDISABLE,
  RXDLYALIGNMONENB,	      
  RXDLYALIGNOVERRIDE,
  RXDLYALIGNRESET,
  RXDLYALIGNSWPPRECURB,
  RXDLYALIGNUPDSW,
  RXENCHANSYNC,
  RXENMCOMMAALIGN,
  RXENPCOMMAALIGN,
  RXENPMAPHASEALIGN,
  RXENPRBSTST,
  RXENSAMPLEALIGN,
  RXEQMIX,
  RXGEARBOXSLIP,
  RXN,
  RXP,
  RXPLLLKDETEN,
  RXPLLPOWERDOWN,
  RXPLLREFSELDY,
  RXPMASETPHASE,
  RXPOLARITY,
  RXPOWERDOWN,
  RXRATE,
  RXRESET,
  RXSLIDE,
  RXUSRCLK,
  RXUSRCLK2,
  SOUTHREFCLKRX,
  SOUTHREFCLKTX,
  TSTCLK0,
  TSTCLK1,
  TSTIN,
  TXBUFDIFFCTRL,
  TXBYPASS8B10B,
  TXCHARDISPMODE,
  TXCHARDISPVAL,
  TXCHARISK,
  TXCOMINIT,
  TXCOMSAS,
  TXCOMWAKE,
  TXDATA,
  TXDEEMPH,
  TXDETECTRX,
  TXDIFFCTRL,
  TXDLYALIGNDISABLE,
  TXDLYALIGNMONENB,    
  TXDLYALIGNOVERRIDE,
  TXDLYALIGNRESET,
  TXDLYALIGNUPDSW,
  TXELECIDLE,
  TXENC8B10BUSE,
  TXENPMAPHASEALIGN,
  TXENPRBSTST,
  TXHEADER,
  TXINHIBIT,
  TXMARGIN,
  TXPDOWNASYNCH,
  TXPLLLKDETEN,
  TXPLLPOWERDOWN,
  TXPLLREFSELDY,
  TXPMASETPHASE,
  TXPOLARITY,
  TXPOSTEMPHASIS,
  TXPOWERDOWN,
  TXPRBSFORCEERR,
  TXPREEMPHASIS,
  TXRATE,
  TXRESET,
  TXSEQUENCE,
  TXSTARTSEQ,
  TXSWING,
  TXUSRCLK,
  TXUSRCLK2,
  USRCODEERR
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input DCLK ;
input DEN ;
input DFEDLYOVRD ;
input DFETAPOVRD ;
input DWE ;
input GATERXELECIDLE ;
input GREFCLKRX ;
input GREFCLKTX ;
input GTXRXRESET ;
input GTXTXRESET ;
input IGNORESIGDET ;
input PERFCLKRX ;
input PERFCLKTX ;
input PLLRXRESET ;
input PLLTXRESET ;
input PRBSCNTRESET ;
input RXBUFRESET ;
input RXCDRRESET ;
input RXCHBONDMASTER ;
input RXCHBONDSLAVE ;
input RXCOMMADETUSE ;
input RXDEC8B10BUSE ;
input RXDLYALIGNDISABLE ;
input RXDLYALIGNMONENB ;
input RXDLYALIGNOVERRIDE ;
input RXDLYALIGNRESET ;
input RXDLYALIGNSWPPRECURB ;
input RXDLYALIGNUPDSW ;
input RXENCHANSYNC ;
input RXENMCOMMAALIGN ;
input RXENPCOMMAALIGN ;
input RXENPMAPHASEALIGN ;
input RXENSAMPLEALIGN ;
input RXGEARBOXSLIP ;
input RXN ;
input RXP ;
input RXPLLLKDETEN ;
input RXPLLPOWERDOWN ;
input RXPMASETPHASE ;
input RXPOLARITY ;
input RXRESET ;
input RXSLIDE ;
input RXUSRCLK2 ;
input RXUSRCLK ;
input TSTCLK0 ;
input TSTCLK1 ;
input TXCOMINIT ;
input TXCOMSAS ;
input TXCOMWAKE ;
input TXDEEMPH ;
input TXDETECTRX ;
input TXDLYALIGNDISABLE ;
input TXDLYALIGNMONENB ;
input TXDLYALIGNOVERRIDE ;
input TXDLYALIGNRESET ;
input TXDLYALIGNUPDSW ;
input TXELECIDLE ;
input TXENC8B10BUSE ;
input TXENPMAPHASEALIGN ;
input TXINHIBIT ;
input TXPDOWNASYNCH ;
input TXPLLLKDETEN ;
input TXPLLPOWERDOWN ;
input TXPMASETPHASE ;
input TXPOLARITY ;
input TXPRBSFORCEERR ;
input TXRESET ;
input TXSTARTSEQ ;
input TXSWING ;
input TXUSRCLK2 ;
input TXUSRCLK ;
input USRCODEERR ;
input [12:0] GTXTEST ;
input [15:0] DI ;
input [19:0] TSTIN ;
input [1:0] MGTREFCLKRX ;
input [1:0] MGTREFCLKTX ;
input [1:0] NORTHREFCLKRX ;
input [1:0] NORTHREFCLKTX ;
input [1:0] RXPOWERDOWN ;
input [1:0] RXRATE ;
input [1:0] SOUTHREFCLKRX ;
input [1:0] SOUTHREFCLKTX ;
input [1:0] TXPOWERDOWN ;
input [1:0] TXRATE ;
input [2:0] LOOPBACK ;
input [2:0] RXCHBONDLEVEL ;
input [2:0] RXENPRBSTST ;
input [2:0] RXPLLREFSELDY ;
input [2:0] TXBUFDIFFCTRL ;
input [2:0] TXENPRBSTST ;
input [2:0] TXHEADER ;
input [2:0] TXMARGIN ;
input [2:0] TXPLLREFSELDY ;
input [31:0] TXDATA ;
input [3:0] DFETAP3 ;
input [3:0] DFETAP4 ;
input [3:0] RXCHBONDI ;
input [3:0] TXBYPASS8B10B ;
input [3:0] TXCHARDISPMODE ;
input [3:0] TXCHARDISPVAL ;
input [3:0] TXCHARISK ;
input [3:0] TXDIFFCTRL ;
input [3:0] TXPREEMPHASIS ;
input [4:0] DFETAP1 ;
input [4:0] DFETAP2 ;
input [4:0] TXPOSTEMPHASIS ;
input [5:0] DFECLKDLYADJ ;
input [6:0] TXSEQUENCE ;
input [7:0] DADDR ;
input [9:0] RXEQMIX ;
output COMFINISH ;
output COMINITDET ;
output COMSASDET ;
output COMWAKEDET ;
output DRDY ;
output PHYSTATUS ;
output RXBYTEISALIGNED ;
output RXBYTEREALIGN ;
output RXCHANBONDSEQ ;
output RXCHANISALIGNED ;
output RXCHANREALIGN ;
output RXCOMMADET ;
output RXDATAVALID ;
output RXELECIDLE ;
output RXHEADERVALID ;
output RXOVERSAMPLEERR ;
output RXPLLLKDET ;
output RXPRBSERR ;
output RXRATEDONE ;
output RXRECCLK ;
output RXRECCLKPCS ;
output RXRESETDONE ;
output RXSTARTOFSEQ ;
output RXVALID ;
output TXGEARBOXREADY ;
output TXN ;
output TXOUTCLK ;
output TXOUTCLKPCS ;
output TXP ;
output TXPLLLKDET ;
output TXRATEDONE ;
output TXRESETDONE ;
output [15:0] DRPDO ;
output [1:0] MGTREFCLKFAB ;
output [1:0] RXLOSSOFSYNC ;
output [1:0] TXBUFSTATUS ;
output [2:0] DFESENSCAL ;
output [2:0] RXBUFSTATUS ;
output [2:0] RXCLKCORCNT ;
output [2:0] RXHEADER ;
output [2:0] RXSTATUS ;
output [31:0] RXDATA ;
output [3:0] DFETAP3MONITOR ;
output [3:0] DFETAP4MONITOR ;
output [3:0] RXCHARISCOMMA ;
output [3:0] RXCHARISK ;
output [3:0] RXCHBONDO ;
output [3:0] RXDISPERR ;
output [3:0] RXNOTINTABLE ;
output [3:0] RXRUNDISP ;
output [3:0] TXKERR ;
output [3:0] TXRUNDISP ;
output [4:0] DFEEYEDACMON ;
output [4:0] DFETAP1MONITOR ;
output [4:0] DFETAP2MONITOR ;
output [5:0] DFECLKDLYADJMON ;
output [7:0] RXDLYALIGNMONITOR ;
output [7:0] TXDLYALIGNMONITOR ;
output [9:0] TSTOUT ;
parameter AC_CAP_DIS = "TRUE";
parameter ALIGN_COMMA_WORD = 1;
parameter [1:0] BGTEST_CFG = 2'b00;
parameter [16:0] BIAS_CFG = 17'h00000;
parameter [4:0] CDR_PH_ADJ_TIME = 5'b10100;
parameter CHAN_BOND_1_MAX_SKEW = 7;
parameter CHAN_BOND_2_MAX_SKEW = 1;
parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0110111100;
parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0110111100;
parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100111100;
parameter [4:0] CHAN_BOND_SEQ_2_CFG = 5'b00000;
parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
parameter CHAN_BOND_SEQ_2_USE = "FALSE";
parameter CHAN_BOND_SEQ_LEN = 1;
parameter CLK_CORRECT_USE = "TRUE";
parameter CLK_COR_ADJ_LEN = 1;
parameter CLK_COR_DET_LEN = 1;
parameter CLK_COR_INSERT_IDLE_FLAG = "FALSE";
parameter CLK_COR_KEEP_IDLE = "FALSE";
parameter CLK_COR_MAX_LAT = 20;
parameter CLK_COR_MIN_LAT = 18;
parameter CLK_COR_PRECEDENCE = "TRUE";
parameter CLK_COR_REPEAT_WAIT = 0;
parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0000000000;
parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
parameter CLK_COR_SEQ_2_USE = "FALSE";
parameter [1:0] CM_TRIM = 2'b01;
parameter [9:0] COMMA_10B_ENABLE = 10'b1111111111;
parameter COMMA_DOUBLE = "FALSE";
parameter [3:0] COM_BURST_VAL = 4'b1111;
parameter DEC_MCOMMA_DETECT = "TRUE";
parameter DEC_PCOMMA_DETECT = "TRUE";
parameter DEC_VALID_COMMA_ONLY = "TRUE";
parameter [4:0] DFE_CAL_TIME = 5'b01100;
parameter [7:0] DFE_CFG = 8'b00011011;
parameter [2:0] GEARBOX_ENDEC = 3'b000;
parameter GEN_RXUSRCLK = "TRUE";
parameter GEN_TXUSRCLK = "TRUE";
parameter GTX_CFG_PWRUP = "TRUE";
parameter [9:0] MCOMMA_10B_VALUE = 10'b1010000011;
parameter MCOMMA_DETECT = "TRUE";
parameter [2:0] OOBDETECT_THRESHOLD = 3'b011;
parameter PCI_EXPRESS_MODE = "FALSE";
parameter [9:0] PCOMMA_10B_VALUE = 10'b0101111100;
parameter PCOMMA_DETECT = "TRUE";
parameter PMA_CAS_CLK_EN = "FALSE";
parameter [26:0] PMA_CDR_SCAN = 27'h640404C;
parameter [75:0] PMA_CFG = 76'h0040000040000000003;
parameter [6:0] PMA_RXSYNC_CFG = 7'h00;
parameter [24:0] PMA_RX_CFG = 25'h05CE048;
parameter [19:0] PMA_TX_CFG = 20'h00082;
parameter [9:0] POWER_SAVE = 10'b0000110100;
parameter RCV_TERM_GND = "FALSE";
parameter RCV_TERM_VTTRX = "TRUE";
parameter RXGEARBOX_USE = "FALSE";
parameter [23:0] RXPLL_COM_CFG = 24'h21680A;
parameter [7:0] RXPLL_CP_CFG = 8'h00;
parameter RXPLL_DIVSEL45_FB = 5;
parameter RXPLL_DIVSEL_FB = 2;
parameter RXPLL_DIVSEL_OUT = 1;
parameter RXPLL_DIVSEL_REF = 1;
parameter [2:0] RXPLL_LKDET_CFG = 3'b111;
parameter [0:0] RXPRBSERR_LOOPBACK = 1'b0;
parameter RXRECCLK_CTRL = "RXRECCLKPCS";
parameter [9:0] RXRECCLK_DLY = 10'b0000000000;
parameter [15:0] RXUSRCLK_DLY = 16'h0000;
parameter RX_BUFFER_USE = "TRUE";
parameter RX_CLK25_DIVIDER = 6;
parameter RX_DATA_WIDTH = 20;
parameter RX_DECODE_SEQ_MATCH = "TRUE";
parameter [3:0] RX_DLYALIGN_CTRINC = 4'b0100;
parameter [4:0] RX_DLYALIGN_EDGESET = 5'b00110;
parameter [3:0] RX_DLYALIGN_LPFINC = 4'b0111;
parameter [2:0] RX_DLYALIGN_MONSEL = 3'b000;
parameter [7:0] RX_DLYALIGN_OVRDSETTING = 8'b00000000;
parameter RX_EN_IDLE_HOLD_CDR = "FALSE";
parameter RX_EN_IDLE_HOLD_DFE = "TRUE";
parameter RX_EN_IDLE_RESET_BUF = "TRUE";
parameter RX_EN_IDLE_RESET_FR = "TRUE";
parameter RX_EN_IDLE_RESET_PH = "TRUE";
parameter RX_EN_MODE_RESET_BUF = "TRUE";
parameter RX_EN_RATE_RESET_BUF = "TRUE";
parameter RX_EN_REALIGN_RESET_BUF = "FALSE";
parameter RX_EN_REALIGN_RESET_BUF2 = "FALSE";
parameter [7:0] RX_EYE_OFFSET = 8'h4C;
parameter [1:0] RX_EYE_SCANMODE = 2'b00;
parameter RX_FIFO_ADDR_MODE = "FULL";
parameter [3:0] RX_IDLE_HI_CNT = 4'b1000;
parameter [3:0] RX_IDLE_LO_CNT = 4'b0000;
parameter RX_LOSS_OF_SYNC_FSM = "FALSE";
parameter RX_LOS_INVALID_INCR = 1;
parameter RX_LOS_THRESHOLD = 4;
parameter RX_OVERSAMPLE_MODE = "FALSE";
parameter RX_SLIDE_AUTO_WAIT = 5;
parameter RX_SLIDE_MODE = "OFF";
parameter RX_XCLK_SEL = "RXREC";
parameter SAS_MAX_COMSAS = 52;
parameter SAS_MIN_COMSAS = 40;
parameter [2:0] SATA_BURST_VAL = 3'b100;
parameter [2:0] SATA_IDLE_VAL = 3'b100;
parameter SATA_MAX_BURST = 7;
parameter SATA_MAX_INIT = 22;
parameter SATA_MAX_WAKE = 7;
parameter SATA_MIN_BURST = 4;
parameter SATA_MIN_INIT = 12;
parameter SATA_MIN_WAKE = 4;
parameter SHOW_REALIGN_COMMA = "TRUE";
parameter SIM_GTXRESET_SPEEDUP = 1;
parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
parameter [2:0] SIM_RXREFCLK_SOURCE = 3'b000;
parameter [2:0] SIM_TXREFCLK_SOURCE = 3'b000;
parameter SIM_TX_ELEC_IDLE_LEVEL = "X";
parameter SIM_VERSION = "2.0";
parameter [4:0] TERMINATION_CTRL = 5'b10100;
parameter TERMINATION_OVRD = "FALSE";
parameter [11:0] TRANS_TIME_FROM_P2 = 12'h03C;
parameter [7:0] TRANS_TIME_NON_P2 = 8'h19;
parameter [7:0] TRANS_TIME_RATE = 8'h0E;
parameter [9:0] TRANS_TIME_TO_P2 = 10'h064;
parameter [31:0] TST_ATTR = 32'h00000000;
parameter TXDRIVE_LOOPBACK_HIZ = "FALSE";
parameter TXDRIVE_LOOPBACK_PD = "FALSE";
parameter TXGEARBOX_USE = "FALSE";
parameter TXOUTCLK_CTRL = "TXOUTCLKPCS";
parameter [9:0] TXOUTCLK_DLY = 10'b0000000000;
parameter [23:0] TXPLL_COM_CFG = 24'h21680A;
parameter [7:0] TXPLL_CP_CFG = 8'h00;
parameter TXPLL_DIVSEL45_FB = 5;
parameter TXPLL_DIVSEL_FB = 2;
parameter TXPLL_DIVSEL_OUT = 1;
parameter TXPLL_DIVSEL_REF = 1;
parameter [2:0] TXPLL_LKDET_CFG = 3'b111;
parameter [1:0] TXPLL_SATA = 2'b00;
parameter TX_BUFFER_USE = "TRUE";
parameter [5:0] TX_BYTECLK_CFG = 6'h00;
parameter TX_CLK25_DIVIDER = 6;
parameter TX_CLK_SOURCE = "RXPLL";
parameter TX_DATA_WIDTH = 20;
parameter [4:0] TX_DEEMPH_0 = 5'b11010;
parameter [4:0] TX_DEEMPH_1 = 5'b10000;
parameter [13:0] TX_DETECT_RX_CFG = 14'h1832;
parameter [3:0] TX_DLYALIGN_CTRINC = 4'b0100;
parameter [3:0] TX_DLYALIGN_LPFINC = 4'b0110;
parameter [2:0] TX_DLYALIGN_MONSEL = 3'b000;
parameter [7:0] TX_DLYALIGN_OVRDSETTING = 8'b10000000;
parameter TX_DRIVE_MODE = "DIRECT";
parameter TX_EN_RATE_RESET_BUF = "TRUE";
parameter [2:0] TX_IDLE_ASSERT_DELAY = 3'b100;
parameter [2:0] TX_IDLE_DEASSERT_DELAY = 3'b010;
parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
parameter TX_OVERSAMPLE_MODE = "FALSE";
parameter [0:0] TX_PMADATA_OPT = 1'b0;
parameter [1:0] TX_TDCC_CFG = 2'b11;
parameter [5:0] TX_USRCLK_CFG = 6'h00;
parameter TX_XCLK_SEL = "TXUSR";
endmodule
//#### END MODULE DEFINITION FOR: GTXE1 ####

//#### BEGIN MODULE DEFINITION FOR :GTXE2_CHANNEL ###
module GTXE2_CHANNEL (
  CPLLFBCLKLOST,
  CPLLLOCK,
  CPLLREFCLKLOST,
  DMONITOROUT,
  DRPDO,
  DRPRDY,
  EYESCANDATAERROR,
  GTREFCLKMONITOR,
  GTXTXN,
  GTXTXP,
  PCSRSVDOUT,
  PHYSTATUS,
  RXBUFSTATUS,
  RXBYTEISALIGNED,
  RXBYTEREALIGN,
  RXCDRLOCK,
  RXCHANBONDSEQ,
  RXCHANISALIGNED,
  RXCHANREALIGN,
  RXCHARISCOMMA,
  RXCHARISK,
  RXCHBONDO,
  RXCLKCORCNT,
  RXCOMINITDET,
  RXCOMMADET,
  RXCOMSASDET,
  RXCOMWAKEDET,
  RXDATA,
  RXDATAVALID,
  RXDISPERR,
  RXDLYSRESETDONE,
  RXELECIDLE,
  RXHEADER,
  RXHEADERVALID,
  RXMONITOROUT,
  RXNOTINTABLE,
  RXOUTCLK,
  RXOUTCLKFABRIC,
  RXOUTCLKPCS,
  RXPHALIGNDONE,
  RXPHMONITOR,
  RXPHSLIPMONITOR,
  RXPRBSERR,
  RXQPISENN,
  RXQPISENP,
  RXRATEDONE,
  RXRESETDONE,
  RXSTARTOFSEQ,
  RXSTATUS,
  RXVALID,
  TSTOUT,
  TXBUFSTATUS,
  TXCOMFINISH,
  TXDLYSRESETDONE,
  TXGEARBOXREADY,
  TXOUTCLK,
  TXOUTCLKFABRIC,
  TXOUTCLKPCS,
  TXPHALIGNDONE,
  TXPHINITDONE,
  TXQPISENN,
  TXQPISENP,
  TXRATEDONE,
  TXRESETDONE,

  CFGRESET,
  CLKRSVD,
  CPLLLOCKDETCLK,
  CPLLLOCKEN,
  CPLLPD,
  CPLLREFCLKSEL,
  CPLLRESET,
  DRPADDR,
  DRPCLK,
  DRPDI,
  DRPEN,
  DRPWE,
  EYESCANMODE,
  EYESCANRESET,
  EYESCANTRIGGER,
  GTGREFCLK,
  GTNORTHREFCLK0,
  GTNORTHREFCLK1,
  GTREFCLK0,
  GTREFCLK1,
  GTRESETSEL,
  GTRSVD,
  GTRXRESET,
  GTSOUTHREFCLK0,
  GTSOUTHREFCLK1,
  GTTXRESET,
  GTXRXN,
  GTXRXP,
  LOOPBACK,
  PCSRSVDIN,
  PCSRSVDIN2,
  PMARSVDIN,
  PMARSVDIN2,
  QPLLCLK,
  QPLLREFCLK,
  RESETOVRD,
  RX8B10BEN,
  RXBUFRESET,
  RXCDRFREQRESET,
  RXCDRHOLD,
  RXCDROVRDEN,
  RXCDRRESET,
  RXCDRRESETRSV,
  RXCHBONDEN,
  RXCHBONDI,
  RXCHBONDLEVEL,
  RXCHBONDMASTER,
  RXCHBONDSLAVE,
  RXCOMMADETEN,
  RXDDIEN,
  RXDFEAGCHOLD,
  RXDFEAGCOVRDEN,
  RXDFECM1EN,
  RXDFELFHOLD,
  RXDFELFOVRDEN,
  RXDFELPMRESET,
  RXDFETAP2HOLD,
  RXDFETAP2OVRDEN,
  RXDFETAP3HOLD,
  RXDFETAP3OVRDEN,
  RXDFETAP4HOLD,
  RXDFETAP4OVRDEN,
  RXDFETAP5HOLD,
  RXDFETAP5OVRDEN,
  RXDFEUTHOLD,
  RXDFEUTOVRDEN,
  RXDFEVPHOLD,
  RXDFEVPOVRDEN,
  RXDFEVSEN,
  RXDFEXYDEN,
  RXDFEXYDHOLD,
  RXDFEXYDOVRDEN,
  RXDLYBYPASS,
  RXDLYEN,
  RXDLYOVRDEN,
  RXDLYSRESET,
  RXELECIDLEMODE,
  RXGEARBOXSLIP,
  RXLPMEN,
  RXLPMHFHOLD,
  RXLPMHFOVRDEN,
  RXLPMLFHOLD,
  RXLPMLFKLOVRDEN,
  RXMCOMMAALIGNEN,
  RXMONITORSEL,
  RXOOBRESET,
  RXOSHOLD,
  RXOSOVRDEN,
  RXOUTCLKSEL,
  RXPCOMMAALIGNEN,
  RXPCSRESET,
  RXPD,
  RXPHALIGN,
  RXPHALIGNEN,
  RXPHDLYPD,
  RXPHDLYRESET,
  RXPHOVRDEN,
  RXPMARESET,
  RXPOLARITY,
  RXPRBSCNTRESET,
  RXPRBSSEL,
  RXQPIEN,
  RXRATE,
  RXSLIDE,
  RXSYSCLKSEL,
  RXUSERRDY,
  RXUSRCLK,
  RXUSRCLK2,
  SETERRSTATUS,
  TSTIN,
  TX8B10BBYPASS,
  TX8B10BEN,
  TXBUFDIFFCTRL,
  TXCHARDISPMODE,
  TXCHARDISPVAL,
  TXCHARISK,
  TXCOMINIT,
  TXCOMSAS,
  TXCOMWAKE,
  TXDATA,
  TXDEEMPH,
  TXDETECTRX,
  TXDIFFCTRL,
  TXDIFFPD,
  TXDLYBYPASS,
  TXDLYEN,
  TXDLYHOLD,
  TXDLYOVRDEN,
  TXDLYSRESET,
  TXDLYUPDOWN,
  TXELECIDLE,
  TXHEADER,
  TXINHIBIT,
  TXMAINCURSOR,
  TXMARGIN,
  TXOUTCLKSEL,
  TXPCSRESET,
  TXPD,
  TXPDELECIDLEMODE,
  TXPHALIGN,
  TXPHALIGNEN,
  TXPHDLYPD,
  TXPHDLYRESET,
  TXPHDLYTSTCLK,
  TXPHINIT,
  TXPHOVRDEN,
  TXPISOPD,
  TXPMARESET,
  TXPOLARITY,
  TXPOSTCURSOR,
  TXPOSTCURSORINV,
  TXPRBSFORCEERR,
  TXPRBSSEL,
  TXPRECURSOR,
  TXPRECURSORINV,
  TXQPIBIASEN,
  TXQPISTRONGPDOWN,
  TXQPIWEAKPUP,
  TXRATE,
  TXSEQUENCE,
  TXSTARTSEQ,
  TXSWING,
  TXSYSCLKSEL,
  TXUSERRDY,
  TXUSRCLK,
  TXUSRCLK2
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CFGRESET ;
input CPLLLOCKDETCLK ;
input CPLLLOCKEN ;
input CPLLPD ;
input CPLLRESET ;
input DRPCLK ;
input DRPEN ;
input DRPWE ;
input EYESCANMODE ;
input EYESCANRESET ;
input EYESCANTRIGGER ;
input GTGREFCLK ;
input GTNORTHREFCLK0 ;
input GTNORTHREFCLK1 ;
input GTREFCLK0 ;
input GTREFCLK1 ;
input GTRESETSEL ;
input GTRXRESET ;
input GTSOUTHREFCLK0 ;
input GTSOUTHREFCLK1 ;
input GTTXRESET ;
input GTXRXN ;
input GTXRXP ;
input QPLLCLK ;
input QPLLREFCLK ;
input RESETOVRD ;
input RX8B10BEN ;
input RXBUFRESET ;
input RXCDRFREQRESET ;
input RXCDRHOLD ;
input RXCDROVRDEN ;
input RXCDRRESET ;
input RXCDRRESETRSV ;
input RXCHBONDEN ;
input RXCHBONDMASTER ;
input RXCHBONDSLAVE ;
input RXCOMMADETEN ;
input RXDDIEN ;
input RXDFEAGCHOLD ;
input RXDFEAGCOVRDEN ;
input RXDFECM1EN ;
input RXDFELFHOLD ;
input RXDFELFOVRDEN ;
input RXDFELPMRESET ;
input RXDFETAP2HOLD ;
input RXDFETAP2OVRDEN ;
input RXDFETAP3HOLD ;
input RXDFETAP3OVRDEN ;
input RXDFETAP4HOLD ;
input RXDFETAP4OVRDEN ;
input RXDFETAP5HOLD ;
input RXDFETAP5OVRDEN ;
input RXDFEUTHOLD ;
input RXDFEUTOVRDEN ;
input RXDFEVPHOLD ;
input RXDFEVPOVRDEN ;
input RXDFEVSEN ;
input RXDFEXYDEN ;
input RXDFEXYDHOLD ;
input RXDFEXYDOVRDEN ;
input RXDLYBYPASS ;
input RXDLYEN ;
input RXDLYOVRDEN ;
input RXDLYSRESET ;
input RXGEARBOXSLIP ;
input RXLPMEN ;
input RXLPMHFHOLD ;
input RXLPMHFOVRDEN ;
input RXLPMLFHOLD ;
input RXLPMLFKLOVRDEN ;
input RXMCOMMAALIGNEN ;
input RXOOBRESET ;
input RXOSHOLD ;
input RXOSOVRDEN ;
input RXPCOMMAALIGNEN ;
input RXPCSRESET ;
input RXPHALIGN ;
input RXPHALIGNEN ;
input RXPHDLYPD ;
input RXPHDLYRESET ;
input RXPHOVRDEN ;
input RXPMARESET ;
input RXPOLARITY ;
input RXPRBSCNTRESET ;
input RXQPIEN ;
input RXSLIDE ;
input RXUSERRDY ;
input RXUSRCLK2 ;
input RXUSRCLK ;
input SETERRSTATUS ;
input TX8B10BEN ;
input TXCOMINIT ;
input TXCOMSAS ;
input TXCOMWAKE ;
input TXDEEMPH ;
input TXDETECTRX ;
input TXDIFFPD ;
input TXDLYBYPASS ;
input TXDLYEN ;
input TXDLYHOLD ;
input TXDLYOVRDEN ;
input TXDLYSRESET ;
input TXDLYUPDOWN ;
input TXELECIDLE ;
input TXINHIBIT ;
input TXPCSRESET ;
input TXPDELECIDLEMODE ;
input TXPHALIGN ;
input TXPHALIGNEN ;
input TXPHDLYPD ;
input TXPHDLYRESET ;
input TXPHDLYTSTCLK ;
input TXPHINIT ;
input TXPHOVRDEN ;
input TXPISOPD ;
input TXPMARESET ;
input TXPOLARITY ;
input TXPOSTCURSORINV ;
input TXPRBSFORCEERR ;
input TXPRECURSORINV ;
input TXQPIBIASEN ;
input TXQPISTRONGPDOWN ;
input TXQPIWEAKPUP ;
input TXSTARTSEQ ;
input TXSWING ;
input TXUSERRDY ;
input TXUSRCLK2 ;
input TXUSRCLK ;
input [15:0] DRPDI ;
input [15:0] GTRSVD ;
input [15:0] PCSRSVDIN ;
input [19:0] TSTIN ;
input [1:0] RXELECIDLEMODE ;
input [1:0] RXMONITORSEL ;
input [1:0] RXPD ;
input [1:0] RXSYSCLKSEL ;
input [1:0] TXPD ;
input [1:0] TXSYSCLKSEL ;
input [2:0] CPLLREFCLKSEL ;
input [2:0] LOOPBACK ;
input [2:0] RXCHBONDLEVEL ;
input [2:0] RXOUTCLKSEL ;
input [2:0] RXPRBSSEL ;
input [2:0] RXRATE ;
input [2:0] TXBUFDIFFCTRL ;
input [2:0] TXHEADER ;
input [2:0] TXMARGIN ;
input [2:0] TXOUTCLKSEL ;
input [2:0] TXPRBSSEL ;
input [2:0] TXRATE ;
input [3:0] CLKRSVD ;
input [3:0] TXDIFFCTRL ;
input [4:0] PCSRSVDIN2 ;
input [4:0] PMARSVDIN2 ;
input [4:0] PMARSVDIN ;
input [4:0] RXCHBONDI ;
input [4:0] TXPOSTCURSOR ;
input [4:0] TXPRECURSOR ;
input [63:0] TXDATA ;
input [6:0] TXMAINCURSOR ;
input [6:0] TXSEQUENCE ;
input [7:0] TX8B10BBYPASS ;
input [7:0] TXCHARDISPMODE ;
input [7:0] TXCHARDISPVAL ;
input [7:0] TXCHARISK ;
input [8:0] DRPADDR ;
output CPLLFBCLKLOST ;
output CPLLLOCK ;
output CPLLREFCLKLOST ;
output DRPRDY ;
output EYESCANDATAERROR ;
output GTREFCLKMONITOR ;
output GTXTXN ;
output GTXTXP ;
output PHYSTATUS ;
output RXBYTEISALIGNED ;
output RXBYTEREALIGN ;
output RXCDRLOCK ;
output RXCHANBONDSEQ ;
output RXCHANISALIGNED ;
output RXCHANREALIGN ;
output RXCOMINITDET ;
output RXCOMMADET ;
output RXCOMSASDET ;
output RXCOMWAKEDET ;
output RXDATAVALID ;
output RXDLYSRESETDONE ;
output RXELECIDLE ;
output RXHEADERVALID ;
output RXOUTCLK ;
output RXOUTCLKFABRIC ;
output RXOUTCLKPCS ;
output RXPHALIGNDONE ;
output RXPRBSERR ;
output RXQPISENN ;
output RXQPISENP ;
output RXRATEDONE ;
output RXRESETDONE ;
output RXSTARTOFSEQ ;
output RXVALID ;
output TXCOMFINISH ;
output TXDLYSRESETDONE ;
output TXGEARBOXREADY ;
output TXOUTCLK ;
output TXOUTCLKFABRIC ;
output TXOUTCLKPCS ;
output TXPHALIGNDONE ;
output TXPHINITDONE ;
output TXQPISENN ;
output TXQPISENP ;
output TXRATEDONE ;
output TXRESETDONE ;
output [15:0] DRPDO ;
output [15:0] PCSRSVDOUT ;
output [1:0] RXCLKCORCNT ;
output [1:0] TXBUFSTATUS ;
output [2:0] RXBUFSTATUS ;
output [2:0] RXHEADER ;
output [2:0] RXSTATUS ;
output [4:0] RXCHBONDO ;
output [4:0] RXPHMONITOR ;
output [4:0] RXPHSLIPMONITOR ;
output [63:0] RXDATA ;
output [6:0] RXMONITOROUT ;
output [7:0] DMONITOROUT ;
output [7:0] RXCHARISCOMMA ;
output [7:0] RXCHARISK ;
output [7:0] RXDISPERR ;
output [7:0] RXNOTINTABLE ;
output [9:0] TSTOUT ;
parameter ALIGN_COMMA_DOUBLE = "FALSE";
parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
parameter ALIGN_COMMA_WORD = 1;
parameter ALIGN_MCOMMA_DET = "TRUE";
parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
parameter ALIGN_PCOMMA_DET = "TRUE";
parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
parameter CBCC_DATA_SOURCE_SEL = "DECODED";
parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
parameter CHAN_BOND_MAX_SKEW = 7;
parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
parameter CHAN_BOND_SEQ_2_USE = "FALSE";
parameter CHAN_BOND_SEQ_LEN = 1;
parameter CLK_CORRECT_USE = "TRUE";
parameter CLK_COR_KEEP_IDLE = "FALSE";
parameter CLK_COR_MAX_LAT = 20;
parameter CLK_COR_MIN_LAT = 18;
parameter CLK_COR_PRECEDENCE = "TRUE";
parameter CLK_COR_REPEAT_WAIT = 0;
parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
parameter CLK_COR_SEQ_2_USE = "FALSE";
parameter CLK_COR_SEQ_LEN = 1;
parameter [23:0] CPLL_CFG = 24'hB007D8;
parameter CPLL_FBDIV = 4;
parameter CPLL_FBDIV_45 = 5;
parameter [23:0] CPLL_INIT_CFG = 24'h00001E;
parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
parameter CPLL_REFCLK_DIV = 1;
parameter DEC_MCOMMA_DETECT = "TRUE";
parameter DEC_PCOMMA_DETECT = "TRUE";
parameter DEC_VALID_COMMA_ONLY = "TRUE";
parameter [23:0] DMONITOR_CFG = 24'h000A00;
parameter [5:0] ES_CONTROL = 6'b000000;
parameter ES_ERRDET_EN = "FALSE";
parameter ES_EYE_SCAN_EN = "FALSE";
parameter [11:0] ES_HORZ_OFFSET = 12'h000;
parameter [9:0] ES_PMA_CFG = 10'b0000000000;
parameter [4:0] ES_PRESCALE = 5'b00000;
parameter [79:0] ES_QUALIFIER = 80'h00000000000000000000;
parameter [79:0] ES_QUAL_MASK = 80'h00000000000000000000;
parameter [79:0] ES_SDATA_MASK = 80'h00000000000000000000;
parameter [8:0] ES_VERT_OFFSET = 9'b000000000;
parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
parameter FTS_LANE_DESKEW_EN = "FALSE";
parameter [2:0] GEARBOX_MODE = 3'b000;
parameter [1:0] OUTREFCLK_SEL_INV = 2'b11;
parameter PCS_PCIE_EN = "FALSE";
parameter [47:0] PCS_RSVD_ATTR = 48'h000000000000;
parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
parameter [31:0] PMA_RSV = 32'h00000000;
parameter [15:0] PMA_RSV2 = 16'h2050;
parameter [1:0] PMA_RSV3 = 2'b00;
parameter [31:0] PMA_RSV4 = 32'h00000000;
parameter [4:0] RXBUFRESET_TIME = 5'b00001;
parameter RXBUF_ADDR_MODE = "FULL";
parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
parameter RXBUF_EN = "TRUE";
parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
parameter RXBUF_RESET_ON_EIDLE = "FALSE";
parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
parameter RXBUF_THRESH_OVFLW = 61;
parameter RXBUF_THRESH_OVRD = "FALSE";
parameter RXBUF_THRESH_UNDFLW = 4;
parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
parameter [71:0] RXCDR_CFG = 72'h0B000023FF20400020;
parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
parameter [5:0] RXCDR_LOCK_CFG = 6'b010101;
parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
parameter [15:0] RXDLY_CFG = 16'h001F;
parameter [8:0] RXDLY_LCFG = 9'h030;
parameter [15:0] RXDLY_TAP_CFG = 16'h0000;
parameter RXGEARBOX_EN = "FALSE";
parameter [4:0] RXISCANRESET_TIME = 5'b00001;
parameter [13:0] RXLPM_HF_CFG = 14'b00000011110000;
parameter [13:0] RXLPM_LF_CFG = 14'b00000011110000;
parameter [6:0] RXOOB_CFG = 7'b0000110;
parameter RXOUT_DIV = 2;
parameter [4:0] RXPCSRESET_TIME = 5'b00001;
parameter [23:0] RXPHDLY_CFG = 24'h084020;
parameter [23:0] RXPH_CFG = 24'h000000;
parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
parameter [4:0] RXPMARESET_TIME = 5'b00011;
parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
parameter RXSLIDE_AUTO_WAIT = 7;
parameter RXSLIDE_MODE = "OFF";
parameter [11:0] RX_BIAS_CFG = 12'b000000000000;
parameter [5:0] RX_BUFFER_CFG = 6'b000000;
parameter RX_CLK25_DIV = 7;
parameter [0:0] RX_CLKMUX_PD = 1'b1;
parameter [1:0] RX_CM_SEL = 2'b11;
parameter [2:0] RX_CM_TRIM = 3'b100;
parameter RX_DATA_WIDTH = 20;
parameter [5:0] RX_DDI_SEL = 6'b000000;
parameter [11:0] RX_DEBUG_CFG = 12'b000000000000;
parameter RX_DEFER_RESET_BUF_EN = "TRUE";
parameter [22:0] RX_DFE_GAIN_CFG = 23'h180E0F;
parameter [11:0] RX_DFE_H2_CFG = 12'b000111100000;
parameter [11:0] RX_DFE_H3_CFG = 12'b000111100000;
parameter [10:0] RX_DFE_H4_CFG = 11'b00011110000;
parameter [10:0] RX_DFE_H5_CFG = 11'b00011110000;
parameter [12:0] RX_DFE_KL_CFG = 13'b0001111110000;
parameter [31:0] RX_DFE_KL_CFG2 = 32'h3008E56A;
parameter [15:0] RX_DFE_LPM_CFG = 16'h0904;
parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
parameter [16:0] RX_DFE_UT_CFG = 17'b00111111000000000;
parameter [16:0] RX_DFE_VP_CFG = 17'b00011111100000000;
parameter [12:0] RX_DFE_XYD_CFG = 13'b0000000010000;
parameter RX_DISPERR_SEQ_MATCH = "TRUE";
parameter RX_INT_DATAWIDTH = 0;
parameter [12:0] RX_OS_CFG = 13'b0001111110000;
parameter RX_SIG_VALID_DLY = 10;
parameter RX_XCLK_SEL = "RXREC";
parameter SAS_MAX_COM = 64;
parameter SAS_MIN_COM = 36;
parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
parameter [2:0] SATA_BURST_VAL = 3'b100;
parameter SATA_CPLL_CFG = "VCO_3000MHZ";
parameter [2:0] SATA_EIDLE_VAL = 3'b100;
parameter SATA_MAX_BURST = 8;
parameter SATA_MAX_INIT = 21;
parameter SATA_MAX_WAKE = 7;
parameter SATA_MIN_BURST = 4;
parameter SATA_MIN_INIT = 12;
parameter SATA_MIN_WAKE = 4;
parameter SHOW_REALIGN_COMMA = "TRUE";
parameter [2:0] SIM_CPLLREFCLK_SEL = 3'b001;
parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
parameter SIM_RESET_SPEEDUP = "TRUE";
parameter SIM_TX_EIDLE_DRIVE_LEVEL = "X";
parameter SIM_VERSION = "4.0";
parameter [4:0] TERM_RCAL_CFG = 5'b10000;
parameter [0:0] TERM_RCAL_OVRD = 1'b0;
parameter [7:0] TRANS_TIME_RATE = 8'h0E;
parameter [31:0] TST_RSV = 32'h00000000;
parameter TXBUF_EN = "TRUE";
parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
parameter [15:0] TXDLY_CFG = 16'h001F;
parameter [8:0] TXDLY_LCFG = 9'h030;
parameter [15:0] TXDLY_TAP_CFG = 16'h0000;
parameter TXGEARBOX_EN = "FALSE";
parameter TXOUT_DIV = 2;
parameter [4:0] TXPCSRESET_TIME = 5'b00001;
parameter [23:0] TXPHDLY_CFG = 24'h084020;
parameter [15:0] TXPH_CFG = 16'h0780;
parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
parameter [4:0] TXPMARESET_TIME = 5'b00001;
parameter TX_CLK25_DIV = 7;
parameter [0:0] TX_CLKMUX_PD = 1'b1;
parameter TX_DATA_WIDTH = 20;
parameter [4:0] TX_DEEMPH0 = 5'b00000;
parameter [4:0] TX_DEEMPH1 = 5'b00000;
parameter TX_DRIVE_MODE = "DIRECT";
parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
parameter TX_INT_DATAWIDTH = 0;
parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
parameter [0:0] TX_PREDRIVER_MODE = 1'b0;
parameter [0:0] TX_QPI_STATUS_EN = 1'b0;
parameter [13:0] TX_RXDETECT_CFG = 14'h1832;
parameter [2:0] TX_RXDETECT_REF = 3'b100;
parameter TX_XCLK_SEL = "TXUSR";
parameter [0:0] UCODEER_CLR = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: GTXE2_CHANNEL ####

//#### BEGIN MODULE DEFINITION FOR :GTXE2_COMMON ###
module GTXE2_COMMON (
  DRPDO,
  DRPRDY,
  QPLLDMONITOR,
  QPLLFBCLKLOST,
  QPLLLOCK,
  QPLLOUTCLK,
  QPLLOUTREFCLK,
  QPLLREFCLKLOST,
  REFCLKOUTMONITOR,

  BGBYPASSB,
  BGMONITORENB,
  BGPDB,
  BGRCALOVRD,
  DRPADDR,
  DRPCLK,
  DRPDI,
  DRPEN,
  DRPWE,
  GTGREFCLK,
  GTNORTHREFCLK0,
  GTNORTHREFCLK1,
  GTREFCLK0,
  GTREFCLK1,
  GTSOUTHREFCLK0,
  GTSOUTHREFCLK1,
  PMARSVD,
  QPLLLOCKDETCLK,
  QPLLLOCKEN,
  QPLLOUTRESET,
  QPLLPD,
  QPLLREFCLKSEL,
  QPLLRESET,
  QPLLRSVD1,
  QPLLRSVD2,
  RCALENB
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input BGBYPASSB ;
input BGMONITORENB ;
input BGPDB ;
input DRPCLK ;
input DRPEN ;
input DRPWE ;
input GTGREFCLK ;
input GTNORTHREFCLK0 ;
input GTNORTHREFCLK1 ;
input GTREFCLK0 ;
input GTREFCLK1 ;
input GTSOUTHREFCLK0 ;
input GTSOUTHREFCLK1 ;
input QPLLLOCKDETCLK ;
input QPLLLOCKEN ;
input QPLLOUTRESET ;
input QPLLPD ;
input QPLLRESET ;
input RCALENB ;
input [15:0] DRPDI ;
input [15:0] QPLLRSVD1 ;
input [2:0] QPLLREFCLKSEL ;
input [4:0] BGRCALOVRD ;
input [4:0] QPLLRSVD2 ;
input [7:0] DRPADDR ;
input [7:0] PMARSVD ;
output DRPRDY ;
output QPLLFBCLKLOST ;
output QPLLLOCK ;
output QPLLOUTCLK ;
output QPLLOUTREFCLK ;
output QPLLREFCLKLOST ;
output REFCLKOUTMONITOR ;
output [15:0] DRPDO ;
output [7:0] QPLLDMONITOR ;
parameter [63:0] BIAS_CFG = 64'h0000040000001000;
parameter [31:0] COMMON_CFG = 32'h00000000;
parameter [26:0] QPLL_CFG = 27'h0680181;
parameter [3:0] QPLL_CLKOUT_CFG = 4'b0000;
parameter [5:0] QPLL_COARSE_FREQ_OVRD = 6'b010000;
parameter [0:0] QPLL_COARSE_FREQ_OVRD_EN = 1'b0;
parameter [9:0] QPLL_CP = 10'b0000011111;
parameter [0:0] QPLL_CP_MONITOR_EN = 1'b0;
parameter [0:0] QPLL_DMONITOR_SEL = 1'b0;
parameter [9:0] QPLL_FBDIV = 10'b0000000000;
parameter [0:0] QPLL_FBDIV_MONITOR_EN = 1'b0;
parameter [0:0] QPLL_FBDIV_RATIO = 1'b0;
parameter [23:0] QPLL_INIT_CFG = 24'h000006;
parameter [15:0] QPLL_LOCK_CFG = 16'h21E8;
parameter [3:0] QPLL_LPF = 4'b1111;
parameter QPLL_REFCLK_DIV = 2;
parameter [2:0] SIM_QPLLREFCLK_SEL = 3'b001;
parameter SIM_RESET_SPEEDUP = "TRUE";
parameter SIM_VERSION = "4.0";
endmodule
//#### END MODULE DEFINITION FOR: GTXE2_COMMON ####

//#### BEGIN MODULE DEFINITION FOR :GTX_DUAL ###
module GTX_DUAL (
	DFECLKDLYADJMONITOR0,
	DFECLKDLYADJMONITOR1,
	DFEEYEDACMONITOR0,
	DFEEYEDACMONITOR1,
	DFESENSCAL0,
	DFESENSCAL1,
	DFETAP1MONITOR0,
	DFETAP1MONITOR1,
	DFETAP2MONITOR0,
	DFETAP2MONITOR1,
	DFETAP3MONITOR0,
	DFETAP3MONITOR1,
	DFETAP4MONITOR0,
	DFETAP4MONITOR1,
	DO,
	DRDY,
	PHYSTATUS0,
	PHYSTATUS1,
	PLLLKDET,
	REFCLKOUT,
	RESETDONE0,
	RESETDONE1,
	RXBUFSTATUS0,
	RXBUFSTATUS1,
	RXBYTEISALIGNED0,
	RXBYTEISALIGNED1,
	RXBYTEREALIGN0,
	RXBYTEREALIGN1,
	RXCHANBONDSEQ0,
	RXCHANBONDSEQ1,
	RXCHANISALIGNED0,
	RXCHANISALIGNED1,
	RXCHANREALIGN0,
	RXCHANREALIGN1,
	RXCHARISCOMMA0,
	RXCHARISCOMMA1,
	RXCHARISK0,
	RXCHARISK1,
	RXCHBONDO0,
	RXCHBONDO1,
	RXCLKCORCNT0,
	RXCLKCORCNT1,
	RXCOMMADET0,
	RXCOMMADET1,
	RXDATA0,
	RXDATA1,
	RXDATAVALID0,
	RXDATAVALID1,
	RXDISPERR0,
	RXDISPERR1,
	RXELECIDLE0,
	RXELECIDLE1,
	RXHEADER0,
	RXHEADER1,
	RXHEADERVALID0,
	RXHEADERVALID1,
	RXLOSSOFSYNC0,
	RXLOSSOFSYNC1,
	RXNOTINTABLE0,
	RXNOTINTABLE1,
	RXOVERSAMPLEERR0,
	RXOVERSAMPLEERR1,
	RXPRBSERR0,
	RXPRBSERR1,
	RXRECCLK0,
	RXRECCLK1,
	RXRUNDISP0,
	RXRUNDISP1,
	RXSTARTOFSEQ0,
	RXSTARTOFSEQ1,
	RXSTATUS0,
	RXSTATUS1,
	RXVALID0,
	RXVALID1,
	TXBUFSTATUS0,
	TXBUFSTATUS1,
	TXGEARBOXREADY0,
	TXGEARBOXREADY1,
	TXKERR0,
	TXKERR1,
	TXN0,
	TXN1,
	TXOUTCLK0,
	TXOUTCLK1,
	TXP0,
	TXP1,
	TXRUNDISP0,
	TXRUNDISP1,

	CLKIN,
	DADDR,
	DCLK,
	DEN,
	DFECLKDLYADJ0,
	DFECLKDLYADJ1,
	DFETAP10,
	DFETAP11,
	DFETAP20,
	DFETAP21,
	DFETAP30,
	DFETAP31,
	DFETAP40,
	DFETAP41,
	DI,
	DWE,
	GTXRESET,
	GTXTEST,
	INTDATAWIDTH,
	LOOPBACK0,
	LOOPBACK1,
	PLLLKDETEN,
	PLLPOWERDOWN,
	PRBSCNTRESET0,
	PRBSCNTRESET1,
	REFCLKPWRDNB,
	RXBUFRESET0,
	RXBUFRESET1,
	RXCDRRESET0,
	RXCDRRESET1,
	RXCHBONDI0,
	RXCHBONDI1,
	RXCOMMADETUSE0,
	RXCOMMADETUSE1,
	RXDATAWIDTH0,
	RXDATAWIDTH1,
	RXDEC8B10BUSE0,
	RXDEC8B10BUSE1,
	RXENCHANSYNC0,
	RXENCHANSYNC1,
	RXENEQB0,
	RXENEQB1,
	RXENMCOMMAALIGN0,
	RXENMCOMMAALIGN1,
	RXENPCOMMAALIGN0,
	RXENPCOMMAALIGN1,
	RXENPMAPHASEALIGN0,
	RXENPMAPHASEALIGN1,
	RXENPRBSTST0,
	RXENPRBSTST1,
	RXENSAMPLEALIGN0,
	RXENSAMPLEALIGN1,
	RXEQMIX0,
	RXEQMIX1,
	RXEQPOLE0,
	RXEQPOLE1,
	RXGEARBOXSLIP0,
	RXGEARBOXSLIP1,
	RXN0,
	RXN1,
	RXP0,
	RXP1,
	RXPMASETPHASE0,
	RXPMASETPHASE1,
	RXPOLARITY0,
	RXPOLARITY1,
	RXPOWERDOWN0,
	RXPOWERDOWN1,
	RXRESET0,
	RXRESET1,
	RXSLIDE0,
	RXSLIDE1,
	RXUSRCLK0,
	RXUSRCLK1,
	RXUSRCLK20,
	RXUSRCLK21,
	TXBUFDIFFCTRL0,
	TXBUFDIFFCTRL1,
	TXBYPASS8B10B0,
	TXBYPASS8B10B1,
	TXCHARDISPMODE0,
	TXCHARDISPMODE1,
	TXCHARDISPVAL0,
	TXCHARDISPVAL1,
	TXCHARISK0,
	TXCHARISK1,
	TXCOMSTART0,
	TXCOMSTART1,
	TXCOMTYPE0,
	TXCOMTYPE1,
	TXDATA0,
	TXDATA1,
	TXDATAWIDTH0,
	TXDATAWIDTH1,
	TXDETECTRX0,
	TXDETECTRX1,
	TXDIFFCTRL0,
	TXDIFFCTRL1,
	TXELECIDLE0,
	TXELECIDLE1,
	TXENC8B10BUSE0,
	TXENC8B10BUSE1,
	TXENPMAPHASEALIGN0,
	TXENPMAPHASEALIGN1,
	TXENPRBSTST0,
	TXENPRBSTST1,
	TXHEADER0,
	TXHEADER1,
	TXINHIBIT0,
	TXINHIBIT1,
	TXPMASETPHASE0,
	TXPMASETPHASE1,
	TXPOLARITY0,
	TXPOLARITY1,
	TXPOWERDOWN0,
	TXPOWERDOWN1,
	TXPREEMPHASIS0,
	TXPREEMPHASIS1,
	TXRESET0,
	TXRESET1,
	TXSEQUENCE0,
	TXSEQUENCE1,
	TXSTARTSEQ0,
	TXSTARTSEQ1,
	TXUSRCLK0,
	TXUSRCLK1,
	TXUSRCLK20,
	TXUSRCLK21

) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKIN ;
input DCLK ;
input DEN ;
input DWE ;
input GTXRESET ;
input INTDATAWIDTH ;
input PLLLKDETEN ;
input PLLPOWERDOWN ;
input PRBSCNTRESET0 ;
input PRBSCNTRESET1 ;
input REFCLKPWRDNB ;
input RXBUFRESET0 ;
input RXBUFRESET1 ;
input RXCDRRESET0 ;
input RXCDRRESET1 ;
input RXCOMMADETUSE0 ;
input RXCOMMADETUSE1 ;
input RXDEC8B10BUSE0 ;
input RXDEC8B10BUSE1 ;
input RXENCHANSYNC0 ;
input RXENCHANSYNC1 ;
input RXENEQB0 ;
input RXENEQB1 ;
input RXENMCOMMAALIGN0 ;
input RXENMCOMMAALIGN1 ;
input RXENPCOMMAALIGN0 ;
input RXENPCOMMAALIGN1 ;
input RXENPMAPHASEALIGN0 ;
input RXENPMAPHASEALIGN1 ;
input RXENSAMPLEALIGN0 ;
input RXENSAMPLEALIGN1 ;
input RXGEARBOXSLIP0 ;
input RXGEARBOXSLIP1 ;
input RXN0 ;
input RXN1 ;
input RXP0 ;
input RXP1 ;
input RXPMASETPHASE0 ;
input RXPMASETPHASE1 ;
input RXPOLARITY0 ;
input RXPOLARITY1 ;
input RXRESET0 ;
input RXRESET1 ;
input RXSLIDE0 ;
input RXSLIDE1 ;
input RXUSRCLK0 ;
input RXUSRCLK1 ;
input RXUSRCLK20 ;
input RXUSRCLK21 ;
input TXCOMSTART0 ;
input TXCOMSTART1 ;
input TXCOMTYPE0 ;
input TXCOMTYPE1 ;
input TXDETECTRX0 ;
input TXDETECTRX1 ;
input TXELECIDLE0 ;
input TXELECIDLE1 ;
input TXENC8B10BUSE0 ;
input TXENC8B10BUSE1 ;
input TXENPMAPHASEALIGN0 ;
input TXENPMAPHASEALIGN1 ;
input TXINHIBIT0 ;
input TXINHIBIT1 ;
input TXPMASETPHASE0 ;
input TXPMASETPHASE1 ;
input TXPOLARITY0 ;
input TXPOLARITY1 ;
input TXRESET0 ;
input TXRESET1 ;
input TXSTARTSEQ0 ;
input TXSTARTSEQ1 ;
input TXUSRCLK0 ;
input TXUSRCLK1 ;
input TXUSRCLK20 ;
input TXUSRCLK21 ;
input [13:0] GTXTEST ;
input [15:0] DI ;
input [1:0] RXDATAWIDTH0 ;
input [1:0] RXDATAWIDTH1 ;
input [1:0] RXENPRBSTST0 ;
input [1:0] RXENPRBSTST1 ;
input [1:0] RXEQMIX0 ;
input [1:0] RXEQMIX1 ;
input [1:0] RXPOWERDOWN0 ;
input [1:0] RXPOWERDOWN1 ;
input [1:0] TXDATAWIDTH0 ;
input [1:0] TXDATAWIDTH1 ;
input [1:0] TXENPRBSTST0 ;
input [1:0] TXENPRBSTST1 ;
input [1:0] TXPOWERDOWN0 ;
input [1:0] TXPOWERDOWN1 ;
input [2:0] LOOPBACK0 ;
input [2:0] LOOPBACK1 ;
input [2:0] TXBUFDIFFCTRL0 ;
input [2:0] TXBUFDIFFCTRL1 ;
input [2:0] TXDIFFCTRL0 ;
input [2:0] TXDIFFCTRL1 ;
input [2:0] TXHEADER0 ;
input [2:0] TXHEADER1 ;
input [31:0] TXDATA0 ;
input [31:0] TXDATA1 ;
input [3:0] DFETAP30 ;
input [3:0] DFETAP31 ;
input [3:0] DFETAP40 ;
input [3:0] DFETAP41 ;
input [3:0] RXCHBONDI0 ;
input [3:0] RXCHBONDI1 ;
input [3:0] RXEQPOLE0 ;
input [3:0] RXEQPOLE1 ;
input [3:0] TXBYPASS8B10B0 ;
input [3:0] TXBYPASS8B10B1 ;
input [3:0] TXCHARDISPMODE0 ;
input [3:0] TXCHARDISPMODE1 ;
input [3:0] TXCHARDISPVAL0 ;
input [3:0] TXCHARDISPVAL1 ;
input [3:0] TXCHARISK0 ;
input [3:0] TXCHARISK1 ;
input [3:0] TXPREEMPHASIS0 ;
input [3:0] TXPREEMPHASIS1 ;
input [4:0] DFETAP10 ;
input [4:0] DFETAP11 ;
input [4:0] DFETAP20 ;
input [4:0] DFETAP21 ;
input [5:0] DFECLKDLYADJ0 ;
input [5:0] DFECLKDLYADJ1 ;
input [6:0] DADDR ;
input [6:0] TXSEQUENCE0 ;
input [6:0] TXSEQUENCE1 ;
output DRDY ;
output PHYSTATUS0 ;
output PHYSTATUS1 ;
output PLLLKDET ;
output REFCLKOUT ;
output RESETDONE0 ;
output RESETDONE1 ;
output RXBYTEISALIGNED0 ;
output RXBYTEISALIGNED1 ;
output RXBYTEREALIGN0 ;
output RXBYTEREALIGN1 ;
output RXCHANBONDSEQ0 ;
output RXCHANBONDSEQ1 ;
output RXCHANISALIGNED0 ;
output RXCHANISALIGNED1 ;
output RXCHANREALIGN0 ;
output RXCHANREALIGN1 ;
output RXCOMMADET0 ;
output RXCOMMADET1 ;
output RXDATAVALID0 ;
output RXDATAVALID1 ;
output RXELECIDLE0 ;
output RXELECIDLE1 ;
output RXHEADERVALID0 ;
output RXHEADERVALID1 ;
output RXOVERSAMPLEERR0 ;
output RXOVERSAMPLEERR1 ;
output RXPRBSERR0 ;
output RXPRBSERR1 ;
output RXRECCLK0 ;
output RXRECCLK1 ;
output RXSTARTOFSEQ0 ;
output RXSTARTOFSEQ1 ;
output RXVALID0 ;
output RXVALID1 ;
output TXGEARBOXREADY0 ;
output TXGEARBOXREADY1 ;
output TXN0 ;
output TXN1 ;
output TXOUTCLK0 ;
output TXOUTCLK1 ;
output TXP0 ;
output TXP1 ;
output [15:0] DO ;
output [1:0] RXLOSSOFSYNC0 ;
output [1:0] RXLOSSOFSYNC1 ;
output [1:0] TXBUFSTATUS0 ;
output [1:0] TXBUFSTATUS1 ;
output [2:0] DFESENSCAL0 ;
output [2:0] DFESENSCAL1 ;
output [2:0] RXBUFSTATUS0 ;
output [2:0] RXBUFSTATUS1 ;
output [2:0] RXCLKCORCNT0 ;
output [2:0] RXCLKCORCNT1 ;
output [2:0] RXHEADER0 ;
output [2:0] RXHEADER1 ;
output [2:0] RXSTATUS0 ;
output [2:0] RXSTATUS1 ;
output [31:0] RXDATA0 ;
output [31:0] RXDATA1 ;
output [3:0] DFETAP3MONITOR0 ;
output [3:0] DFETAP3MONITOR1 ;
output [3:0] DFETAP4MONITOR0 ;
output [3:0] DFETAP4MONITOR1 ;
output [3:0] RXCHARISCOMMA0 ;
output [3:0] RXCHARISCOMMA1 ;
output [3:0] RXCHARISK0 ;
output [3:0] RXCHARISK1 ;
output [3:0] RXCHBONDO0 ;
output [3:0] RXCHBONDO1 ;
output [3:0] RXDISPERR0 ;
output [3:0] RXDISPERR1 ;
output [3:0] RXNOTINTABLE0 ;
output [3:0] RXNOTINTABLE1 ;
output [3:0] RXRUNDISP0 ;
output [3:0] RXRUNDISP1 ;
output [3:0] TXKERR0 ;
output [3:0] TXKERR1 ;
output [3:0] TXRUNDISP0 ;
output [3:0] TXRUNDISP1 ;
output [4:0] DFEEYEDACMONITOR0 ;
output [4:0] DFEEYEDACMONITOR1 ;
output [4:0] DFETAP1MONITOR0 ;
output [4:0] DFETAP1MONITOR1 ;
output [4:0] DFETAP2MONITOR0 ;
output [4:0] DFETAP2MONITOR1 ;
output [5:0] DFECLKDLYADJMONITOR0 ;
output [5:0] DFECLKDLYADJMONITOR1 ;
parameter AC_CAP_DIS_0 = "TRUE";
parameter AC_CAP_DIS_1 = "TRUE";
parameter CHAN_BOND_KEEP_ALIGN_0 = "FALSE";
parameter CHAN_BOND_KEEP_ALIGN_1 = "FALSE";
parameter CHAN_BOND_MODE_0 = "OFF";
parameter CHAN_BOND_MODE_1 = "OFF";
parameter CHAN_BOND_SEQ_2_USE_0 = "FALSE";
parameter CHAN_BOND_SEQ_2_USE_1 = "FALSE";
parameter CLKINDC_B = "TRUE";
parameter CLKRCV_TRST = "TRUE";
parameter CLK_CORRECT_USE_0 = "TRUE";
parameter CLK_CORRECT_USE_1 = "TRUE";
parameter CLK_COR_INSERT_IDLE_FLAG_0 = "FALSE";
parameter CLK_COR_INSERT_IDLE_FLAG_1 = "FALSE";
parameter CLK_COR_KEEP_IDLE_0 = "FALSE";
parameter CLK_COR_KEEP_IDLE_1 = "FALSE";
parameter CLK_COR_PRECEDENCE_0 = "TRUE";
parameter CLK_COR_PRECEDENCE_1 = "TRUE";
parameter CLK_COR_SEQ_2_USE_0 = "FALSE";
parameter CLK_COR_SEQ_2_USE_1 = "FALSE";
parameter COMMA_DOUBLE_0 = "FALSE";
parameter COMMA_DOUBLE_1 = "FALSE";
parameter DEC_MCOMMA_DETECT_0 = "TRUE";
parameter DEC_MCOMMA_DETECT_1 = "TRUE";
parameter DEC_PCOMMA_DETECT_0 = "TRUE";
parameter DEC_PCOMMA_DETECT_1 = "TRUE";
parameter DEC_VALID_COMMA_ONLY_0 = "TRUE";
parameter DEC_VALID_COMMA_ONLY_1 = "TRUE";
parameter MCOMMA_DETECT_0 = "TRUE";
parameter MCOMMA_DETECT_1 = "TRUE";
parameter OVERSAMPLE_MODE = "FALSE";
parameter PCI_EXPRESS_MODE_0 = "FALSE";
parameter PCI_EXPRESS_MODE_1 = "FALSE";
parameter PCOMMA_DETECT_0 = "TRUE";
parameter PCOMMA_DETECT_1 = "TRUE";
parameter PLL_FB_DCCEN = "FALSE";
parameter PLL_SATA_0 = "FALSE";
parameter PLL_SATA_1 = "FALSE";
parameter RCV_TERM_GND_0 = "FALSE";
parameter RCV_TERM_GND_1 = "FALSE";
parameter RCV_TERM_VTTRX_0 = "FALSE";
parameter RCV_TERM_VTTRX_1 = "FALSE";
parameter RXGEARBOX_USE_0 = "FALSE";
parameter RXGEARBOX_USE_1 = "FALSE";
parameter RX_BUFFER_USE_0 = "TRUE";
parameter RX_BUFFER_USE_1 = "TRUE";
parameter RX_DECODE_SEQ_MATCH_0 = "TRUE";
parameter RX_DECODE_SEQ_MATCH_1 = "TRUE";
parameter RX_EN_IDLE_HOLD_CDR = "FALSE";
parameter RX_EN_IDLE_HOLD_DFE_0 = "TRUE";
parameter RX_EN_IDLE_HOLD_DFE_1 = "TRUE";
parameter RX_EN_IDLE_RESET_BUF_0 = "TRUE";
parameter RX_EN_IDLE_RESET_BUF_1 = "TRUE";
parameter RX_EN_IDLE_RESET_FR = "TRUE";
parameter RX_EN_IDLE_RESET_PH = "TRUE";
parameter RX_LOSS_OF_SYNC_FSM_0 = "FALSE";
parameter RX_LOSS_OF_SYNC_FSM_1 = "FALSE";
parameter RX_SLIDE_MODE_0 = "PCS";
parameter RX_SLIDE_MODE_1 = "PCS";
parameter RX_STATUS_FMT_0 = "PCIE";
parameter RX_STATUS_FMT_1 = "PCIE";
parameter RX_XCLK_SEL_0 = "RXREC";
parameter RX_XCLK_SEL_1 = "RXREC";
parameter SIM_MODE = "FAST";
parameter SIM_PLL_PERDIV2 = 9'h140;
parameter SIM_RECEIVER_DETECT_PASS_0 = "TRUE";
parameter SIM_RECEIVER_DETECT_PASS_1 = "TRUE";
parameter TERMINATION_OVRD = "FALSE";
parameter TXGEARBOX_USE_0 = "FALSE";
parameter TXGEARBOX_USE_1 = "FALSE";
parameter TX_BUFFER_USE_0 = "TRUE";
parameter TX_BUFFER_USE_1 = "TRUE";
parameter TX_XCLK_SEL_0 = "TXOUT";
parameter TX_XCLK_SEL_1 = "TXOUT";
parameter [11:0] TRANS_TIME_FROM_P2_0 = 12'h03c;
parameter [11:0] TRANS_TIME_FROM_P2_1 = 12'h03c;
parameter [13:0] TX_DETECT_RX_CFG_0 = 14'h1832;
parameter [13:0] TX_DETECT_RX_CFG_1 = 14'h1832;
parameter [19:0] PMA_TX_CFG_0 = 20'h80082;
parameter [19:0] PMA_TX_CFG_1 = 20'h80082;
parameter [1:0] CM_TRIM_0 = 2'b10;
parameter [1:0] CM_TRIM_1 = 2'b10;
parameter [23:0] PLL_COM_CFG = 24'h21680a;
parameter [24:0] PMA_RX_CFG_0 = 25'h0f44089;
parameter [24:0] PMA_RX_CFG_1 = 25'h0f44089;
parameter [26:0] PMA_CDR_SCAN_0 = 27'h6404035;
parameter [26:0] PMA_CDR_SCAN_1 = 27'h6404035;
parameter [2:0] GEARBOX_ENDEC_0 = 3'b000;
parameter [2:0] GEARBOX_ENDEC_1 = 3'b000;
parameter [2:0] OOBDETECT_THRESHOLD_0 = 3'b110;
parameter [2:0] OOBDETECT_THRESHOLD_1 = 3'b110;
parameter [2:0] PLL_LKDET_CFG = 3'b101;
parameter [2:0] PLL_TDCC_CFG = 3'b000;
parameter [2:0] SATA_BURST_VAL_0 = 3'b100;
parameter [2:0] SATA_BURST_VAL_1 = 3'b100;
parameter [2:0] SATA_IDLE_VAL_0 = 3'b100;
parameter [2:0] SATA_IDLE_VAL_1 = 3'b100;
parameter [2:0] TXRX_INVERT_0 = 3'b011;
parameter [2:0] TXRX_INVERT_1 = 3'b011;
parameter [2:0] TX_IDLE_DELAY_0 = 3'b010;
parameter [2:0] TX_IDLE_DELAY_1 = 3'b010;
parameter [31:0] PRBS_ERR_THRESHOLD_0 = 32'h00000001;
parameter [31:0] PRBS_ERR_THRESHOLD_1 = 32'h00000001;
parameter [3:0] CHAN_BOND_SEQ_1_ENABLE_0 = 4'b0001;
parameter [3:0] CHAN_BOND_SEQ_1_ENABLE_1 = 4'b0001;
parameter [3:0] CHAN_BOND_SEQ_2_ENABLE_0 = 4'b0000;
parameter [3:0] CHAN_BOND_SEQ_2_ENABLE_1 = 4'b0000;
parameter [3:0] CLK_COR_SEQ_1_ENABLE_0 = 4'b0001;
parameter [3:0] CLK_COR_SEQ_1_ENABLE_1 = 4'b0001;
parameter [3:0] CLK_COR_SEQ_2_ENABLE_0 = 4'b0000;
parameter [3:0] CLK_COR_SEQ_2_ENABLE_1 = 4'b0000;
parameter [3:0] COM_BURST_VAL_0 = 4'b1111;
parameter [3:0] COM_BURST_VAL_1 = 4'b1111;
parameter [3:0] RX_IDLE_HI_CNT_0 = 4'b1000;
parameter [3:0] RX_IDLE_HI_CNT_1 = 4'b1000;
parameter [3:0] RX_IDLE_LO_CNT_0 = 4'b0000;
parameter [3:0] RX_IDLE_LO_CNT_1 = 4'b0000;
parameter [4:0] CDR_PH_ADJ_TIME = 5'b01010;
parameter [4:0] DFE_CAL_TIME = 5'b00110;
parameter [4:0] TERMINATION_CTRL = 5'b10100;
parameter [68:0] PMA_COM_CFG = 69'h0;
parameter [6:0] PMA_RXSYNC_CFG_0 = 7'h0;
parameter [6:0] PMA_RXSYNC_CFG_1 = 7'h0;
parameter [7:0] PLL_CP_CFG = 8'h00;
parameter [7:0] TRANS_TIME_NON_P2_0 = 8'h19;
parameter [7:0] TRANS_TIME_NON_P2_1 = 8'h19;
parameter [9:0] CHAN_BOND_SEQ_1_1_0 = 10'b0101111100;
parameter [9:0] CHAN_BOND_SEQ_1_1_1 = 10'b0101111100;
parameter [9:0] CHAN_BOND_SEQ_1_2_0 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_1_2_1 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_1_3_0 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_1_3_1 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_1_4_0 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_1_4_1 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_2_1_0 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_2_1_1 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_2_2_0 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_2_2_1 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_2_3_0 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_2_3_1 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_2_4_0 = 10'b0000000000;
parameter [9:0] CHAN_BOND_SEQ_2_4_1 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_1_0 = 10'b0100011100;
parameter [9:0] CLK_COR_SEQ_1_1_1 = 10'b0100011100;
parameter [9:0] CLK_COR_SEQ_1_2_0 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_2_1 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_3_0 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_3_1 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_4_0 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_1_4_1 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_1_0 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_1_1 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_2_0 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_2_1 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_3_0 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_3_1 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_4_0 = 10'b0000000000;
parameter [9:0] CLK_COR_SEQ_2_4_1 = 10'b0000000000;
parameter [9:0] COMMA_10B_ENABLE_0 = 10'b0001111111;
parameter [9:0] COMMA_10B_ENABLE_1 = 10'b0001111111;
parameter [9:0] DFE_CFG_0 = 10'b1101111011;
parameter [9:0] DFE_CFG_1 = 10'b1101111011;
parameter [9:0] MCOMMA_10B_VALUE_0 = 10'b1010000011;
parameter [9:0] MCOMMA_10B_VALUE_1 = 10'b1010000011;
parameter [9:0] PCOMMA_10B_VALUE_0 = 10'b0101111100;
parameter [9:0] PCOMMA_10B_VALUE_1 = 10'b0101111100;
parameter [9:0] TRANS_TIME_TO_P2_0 = 10'h064;
parameter [9:0] TRANS_TIME_TO_P2_1 = 10'h064;
parameter ALIGN_COMMA_WORD_0 = 1;
parameter ALIGN_COMMA_WORD_1 = 1;
parameter CB2_INH_CC_PERIOD_0 = 8;
parameter CB2_INH_CC_PERIOD_1 = 8;
parameter CHAN_BOND_1_MAX_SKEW_0 = 7;
parameter CHAN_BOND_1_MAX_SKEW_1 = 7;
parameter CHAN_BOND_2_MAX_SKEW_0 = 7;
parameter CHAN_BOND_2_MAX_SKEW_1 = 7;
parameter CHAN_BOND_LEVEL_0 = 0;
parameter CHAN_BOND_LEVEL_1 = 0;
parameter CHAN_BOND_SEQ_LEN_0 = 1;
parameter CHAN_BOND_SEQ_LEN_1 = 1;
parameter CLK25_DIVIDER = 10;
parameter CLK_COR_ADJ_LEN_0 = 1;
parameter CLK_COR_ADJ_LEN_1 = 1;
parameter CLK_COR_DET_LEN_0 = 1;
parameter CLK_COR_DET_LEN_1 = 1;
parameter CLK_COR_MAX_LAT_0 = 20;
parameter CLK_COR_MAX_LAT_1 = 20;
parameter CLK_COR_MIN_LAT_0 = 18;
parameter CLK_COR_MIN_LAT_1 = 18;
parameter CLK_COR_REPEAT_WAIT_0 = 0;
parameter CLK_COR_REPEAT_WAIT_1 = 0;
parameter OOB_CLK_DIVIDER = 6;
parameter PLL_DIVSEL_FB = 2;
parameter PLL_DIVSEL_REF = 1;
parameter PLL_RXDIVSEL_OUT_0 = 1;
parameter PLL_RXDIVSEL_OUT_1 = 1;
parameter PLL_TXDIVSEL_OUT_0 = 1;
parameter PLL_TXDIVSEL_OUT_1 = 1;
parameter RX_LOS_INVALID_INCR_0 = 1;
parameter RX_LOS_INVALID_INCR_1 = 1;
parameter RX_LOS_THRESHOLD_0 = 4;
parameter RX_LOS_THRESHOLD_1 = 4;
parameter SATA_MAX_BURST_0 = 7;
parameter SATA_MAX_BURST_1 = 7;
parameter SATA_MAX_INIT_0 = 22;
parameter SATA_MAX_INIT_1 = 22;
parameter SATA_MAX_WAKE_0 = 7;
parameter SATA_MAX_WAKE_1 = 7;
parameter SATA_MIN_BURST_0 = 4;
parameter SATA_MIN_BURST_1 = 4;
parameter SATA_MIN_INIT_0 = 12;
parameter SATA_MIN_INIT_1 = 12;
parameter SATA_MIN_WAKE_0 = 4;
parameter SATA_MIN_WAKE_1 = 4;
parameter SIM_GTXRESET_SPEEDUP = 1;
parameter TERMINATION_IMP_0 = 50;
parameter TERMINATION_IMP_1 = 50;
endmodule
//#### END MODULE DEFINITION FOR: GTX_DUAL ####

//#### BEGIN MODULE DEFINITION FOR :GTZE2_OCTAL ###
module GTZE2_OCTAL (
  CFGBADVERSIONB,
  CFGCRCERRB,
  CFGGTZDONEB,
  CFGSEUERRB,
  DRPDO,
  DRPRDY,
  DRPSTATUS,
  DRPWDTERR,
  FIBRSVDOUT0,
  FIBRSVDOUT1,
  FIBRSVDOUT2,
  FIBRSVDOUT3,
  FIBRSVDOUT4,
  FIBRSVDOUT5,
  FIBRSVDOUT6,
  FIBRSVDOUT7,
  GTZINITDONEB,
  GTZTXN0,
  GTZTXN1,
  GTZTXN2,
  GTZTXN3,
  GTZTXN4,
  GTZTXN5,
  GTZTXN6,
  GTZTXN7,
  GTZTXP0,
  GTZTXP1,
  GTZTXP2,
  GTZTXP3,
  GTZTXP4,
  GTZTXP5,
  GTZTXP6,
  GTZTXP7,
  RSVDOUT,
  RXDATA0,
  RXDATA1,
  RXDATA2,
  RXDATA3,
  RXDATA4,
  RXDATA5,
  RXDATA6,
  RXDATA7,
  RXDATAVALID0,
  RXDATAVALID1,
  RXDATAVALID2,
  RXDATAVALID3,
  RXDATAVALID4,
  RXDATAVALID5,
  RXDATAVALID6,
  RXDATAVALID7,
  RXFIFOSTATUS0,
  RXFIFOSTATUS1,
  RXFIFOSTATUS2,
  RXFIFOSTATUS3,
  RXFIFOSTATUS4,
  RXFIFOSTATUS5,
  RXFIFOSTATUS6,
  RXFIFOSTATUS7,
  RXHEADER0,
  RXHEADER1,
  RXHEADER2,
  RXHEADER3,
  RXHEADER4,
  RXHEADER5,
  RXHEADER6,
  RXHEADER7,
  RXHEADERVALID0,
  RXHEADERVALID1,
  RXHEADERVALID2,
  RXHEADERVALID3,
  RXHEADERVALID4,
  RXHEADERVALID5,
  RXHEADERVALID6,
  RXHEADERVALID7,
  RXOUTCLK0,
  RXOUTCLK1,
  RXOUTCLK2,
  RXOUTCLK3,
  RXPRBSPASS0,
  RXPRBSPASS1,
  RXPRBSPASS2,
  RXPRBSPASS3,
  RXPRBSPASS4,
  RXPRBSPASS5,
  RXPRBSPASS6,
  RXPRBSPASS7,
  RXRDY0,
  RXRDY1,
  RXRDY2,
  RXRDY3,
  RXRDY4,
  RXRDY5,
  RXRDY6,
  RXRDY7,
  RXRESETDONE0,
  RXRESETDONE1,
  RXRESETDONE2,
  RXRESETDONE3,
  RXRESETDONE4,
  RXRESETDONE5,
  RXRESETDONE6,
  RXRESETDONE7,
  RXSIGNALOK0,
  RXSIGNALOK1,
  RXSIGNALOK2,
  RXSIGNALOK3,
  RXSIGNALOK4,
  RXSIGNALOK5,
  RXSIGNALOK6,
  RXSIGNALOK7,
  SPARESBUSDATAOUT,
  SPARESBUSDONE,
  SPARESBUSRCVDATAVALID,
  SPARESBUSRESULTCODE,
  TXFIFOSTATUS0,
  TXFIFOSTATUS1,
  TXFIFOSTATUS2,
  TXFIFOSTATUS3,
  TXFIFOSTATUS4,
  TXFIFOSTATUS5,
  TXFIFOSTATUS6,
  TXFIFOSTATUS7,
  TXOUTCLK0,
  TXOUTCLK1,
  TXPHASEOUT0,
  TXPHASEOUT1,
  TXPHASEOUT2,
  TXPHASEOUT3,
  TXPHASEOUT4,
  TXPHASEOUT5,
  TXPHASEOUT6,
  TXPHASEOUT7,
  TXRDY0,
  TXRDY1,
  TXRDY2,
  TXRDY3,
  TXRDY4,
  TXRDY5,
  TXRDY6,
  TXRDY7,
  TXRESETDONE0,
  TXRESETDONE1,
  TXRESETDONE2,
  TXRESETDONE3,
  TXRESETDONE4,
  TXRESETDONE5,
  TXRESETDONE6,
  TXRESETDONE7,

  CFGCLK,
  CFGDATA,
  CFGDATAVALID,
  CFGDEBUGMODEB,
  CFGFORCESEUERRB,
  CFGREADBACKB,
  CORECNTL0,
  CORECNTL1,
  CORECNTL2,
  CORECNTL3,
  CORECNTL4,
  CORECNTL5,
  CORECNTL6,
  CORECNTL7,
  DRPADDR,
  DRPCLK0,
  DRPCLK1,
  DRPCLKSEL,
  DRPDI,
  DRPEN,
  DRPWE,
  FARLOOPBACKEN0,
  FARLOOPBACKEN1,
  FARLOOPBACKEN2,
  FARLOOPBACKEN3,
  FARLOOPBACKEN4,
  FARLOOPBACKEN5,
  FARLOOPBACKEN6,
  FARLOOPBACKEN7,
  FIBRSVDIN0,
  FIBRSVDIN1,
  FIBRSVDIN2,
  FIBRSVDIN3,
  FIBRSVDIN4,
  FIBRSVDIN5,
  FIBRSVDIN6,
  FIBRSVDIN7,
  GTREFCLK0N,
  GTREFCLK0P,
  GTREFCLK1N,
  GTREFCLK1P,
  GTZINIT,
  GTZRXN0,
  GTZRXN1,
  GTZRXN2,
  GTZRXN3,
  GTZRXN4,
  GTZRXN5,
  GTZRXN6,
  GTZRXN7,
  GTZRXP0,
  GTZRXP1,
  GTZRXP2,
  GTZRXP3,
  GTZRXP4,
  GTZRXP5,
  GTZRXP6,
  GTZRXP7,
  GTZRXRESET0,
  GTZRXRESET1,
  GTZRXRESET2,
  GTZRXRESET3,
  GTZRXRESET4,
  GTZRXRESET5,
  GTZRXRESET6,
  GTZRXRESET7,
  GTZTXRESET0,
  GTZTXRESET1,
  GTZTXRESET2,
  GTZTXRESET3,
  GTZTXRESET4,
  GTZTXRESET5,
  GTZTXRESET6,
  GTZTXRESET7,
  NEARLOOPBACKEN0,
  NEARLOOPBACKEN1,
  NEARLOOPBACKEN2,
  NEARLOOPBACKEN3,
  NEARLOOPBACKEN4,
  NEARLOOPBACKEN5,
  NEARLOOPBACKEN6,
  NEARLOOPBACKEN7,
  PLLRECALEN0,
  PLLRECALEN1,
  PLLRECALEN2,
  PLLRECALEN3,
  PLLRECALEN4,
  PLLRECALEN5,
  PLLRECALEN6,
  PLLRECALEN7,
  REFCLKSEL0,
  REFCLKSEL1,
  REFCLKSEL2,
  REFCLKSEL3,
  REFCLKSEL4,
  REFCLKSEL5,
  REFCLKSEL6,
  REFCLKSEL7,
  REFSEL0,
  REFSEL1,
  REFSEL2,
  REFSEL3,
  REFSEL4,
  REFSEL5,
  REFSEL6,
  REFSEL7,
  RSVDIN,
  RXBITSLIP0,
  RXBITSLIP1,
  RXBITSLIP2,
  RXBITSLIP3,
  RXBITSLIP4,
  RXBITSLIP5,
  RXBITSLIP6,
  RXBITSLIP7,
  RXDATAWIDTH0,
  RXDATAWIDTH1,
  RXDATAWIDTH2,
  RXDATAWIDTH3,
  RXDATAWIDTH4,
  RXDATAWIDTH5,
  RXDATAWIDTH6,
  RXDATAWIDTH7,
  RXEN0,
  RXEN1,
  RXEN2,
  RXEN3,
  RXEN4,
  RXEN5,
  RXEN6,
  RXEN7,
  RXFIBRESET0,
  RXFIBRESET1,
  RXFIBRESET2,
  RXFIBRESET3,
  RXFIBRESET4,
  RXFIBRESET5,
  RXFIBRESET6,
  RXFIBRESET7,
  RXGEARBOXSLIP0,
  RXGEARBOXSLIP1,
  RXGEARBOXSLIP2,
  RXGEARBOXSLIP3,
  RXGEARBOXSLIP4,
  RXGEARBOXSLIP5,
  RXGEARBOXSLIP6,
  RXGEARBOXSLIP7,
  RXLATCLK,
  RXPOLARITY0,
  RXPOLARITY1,
  RXPOLARITY2,
  RXPOLARITY3,
  RXPOLARITY4,
  RXPOLARITY5,
  RXPOLARITY6,
  RXPOLARITY7,
  RXPRBSEN0,
  RXPRBSEN1,
  RXPRBSEN2,
  RXPRBSEN3,
  RXPRBSEN4,
  RXPRBSEN5,
  RXPRBSEN6,
  RXPRBSEN7,
  RXPRBSSEL0,
  RXPRBSSEL1,
  RXPRBSSEL2,
  RXPRBSSEL3,
  RXPRBSSEL4,
  RXPRBSSEL5,
  RXPRBSSEL6,
  RXPRBSSEL7,
  RXRATESEL0,
  RXRATESEL1,
  RXRATESEL2,
  RXRATESEL3,
  RXRATESEL4,
  RXRATESEL5,
  RXRATESEL6,
  RXRATESEL7,
  RXUSRCLK0,
  RXUSRCLK1,
  RXUSRCLK2,
  RXUSRCLK3,
  RXUSRCLK4,
  RXUSRCLK5,
  RXUSRCLK6,
  RXUSRCLK7,
  SBUSCLKSEL,
  SBUSRESETB,
  SPARESBUSCOMMAND,
  SPARESBUSDATA,
  SPARESBUSDATAADDR,
  SPARESBUSEXECUTEB,
  SPARESBUSRCVDATAVALIDSEL,
  SPARESBUSRECADDR,
  TSTRSVD0,
  TSTRSVD1,
  TSTRSVD2,
  TSTRSVD3,
  TSTRSVD4,
  TXATTNCTRL0,
  TXATTNCTRL1,
  TXATTNCTRL2,
  TXATTNCTRL3,
  TXATTNCTRL4,
  TXATTNCTRL5,
  TXATTNCTRL6,
  TXATTNCTRL7,
  TXDATA0,
  TXDATA1,
  TXDATA2,
  TXDATA3,
  TXDATA4,
  TXDATA5,
  TXDATA6,
  TXDATA7,
  TXDATAWIDTH0,
  TXDATAWIDTH1,
  TXDATAWIDTH2,
  TXDATAWIDTH3,
  TXDATAWIDTH4,
  TXDATAWIDTH5,
  TXDATAWIDTH6,
  TXDATAWIDTH7,
  TXEN0,
  TXEN1,
  TXEN2,
  TXEN3,
  TXEN4,
  TXEN5,
  TXEN6,
  TXEN7,
  TXEQPOSTCTRL0,
  TXEQPOSTCTRL1,
  TXEQPOSTCTRL2,
  TXEQPOSTCTRL3,
  TXEQPOSTCTRL4,
  TXEQPOSTCTRL5,
  TXEQPOSTCTRL6,
  TXEQPOSTCTRL7,
  TXEQPRECTRL0,
  TXEQPRECTRL1,
  TXEQPRECTRL2,
  TXEQPRECTRL3,
  TXEQPRECTRL4,
  TXEQPRECTRL5,
  TXEQPRECTRL6,
  TXEQPRECTRL7,
  TXFIBRESET0,
  TXFIBRESET1,
  TXFIBRESET2,
  TXFIBRESET3,
  TXFIBRESET4,
  TXFIBRESET5,
  TXFIBRESET6,
  TXFIBRESET7,
  TXHEADER0,
  TXHEADER1,
  TXHEADER2,
  TXHEADER3,
  TXHEADER4,
  TXHEADER5,
  TXHEADER6,
  TXHEADER7,
  TXLATCLK,
  TXOUTPUTEN0,
  TXOUTPUTEN1,
  TXOUTPUTEN2,
  TXOUTPUTEN3,
  TXOUTPUTEN4,
  TXOUTPUTEN5,
  TXOUTPUTEN6,
  TXOUTPUTEN7,
  TXOVERRIDEEN0,
  TXOVERRIDEEN1,
  TXOVERRIDEEN2,
  TXOVERRIDEEN3,
  TXOVERRIDEEN4,
  TXOVERRIDEEN5,
  TXOVERRIDEEN6,
  TXOVERRIDEEN7,
  TXOVERRIDEIN0,
  TXOVERRIDEIN1,
  TXOVERRIDEIN2,
  TXOVERRIDEIN3,
  TXOVERRIDEIN4,
  TXOVERRIDEIN5,
  TXOVERRIDEIN6,
  TXOVERRIDEIN7,
  TXPHASECALEN0,
  TXPHASECALEN1,
  TXPHASECALEN2,
  TXPHASECALEN3,
  TXPHASECALEN4,
  TXPHASECALEN5,
  TXPHASECALEN6,
  TXPHASECALEN7,
  TXPHASESLIP0,
  TXPHASESLIP1,
  TXPHASESLIP2,
  TXPHASESLIP3,
  TXPHASESLIP4,
  TXPHASESLIP5,
  TXPHASESLIP6,
  TXPHASESLIP7,
  TXPOLARITY0,
  TXPOLARITY1,
  TXPOLARITY2,
  TXPOLARITY3,
  TXPOLARITY4,
  TXPOLARITY5,
  TXPOLARITY6,
  TXPOLARITY7,
  TXPRBSEN0,
  TXPRBSEN1,
  TXPRBSEN2,
  TXPRBSEN3,
  TXPRBSEN4,
  TXPRBSEN5,
  TXPRBSEN6,
  TXPRBSEN7,
  TXPRBSSEL0,
  TXPRBSSEL1,
  TXPRBSSEL2,
  TXPRBSSEL3,
  TXPRBSSEL4,
  TXPRBSSEL5,
  TXPRBSSEL6,
  TXPRBSSEL7,
  TXRATESEL0,
  TXRATESEL1,
  TXRATESEL2,
  TXRATESEL3,
  TXRATESEL4,
  TXRATESEL5,
  TXRATESEL6,
  TXRATESEL7,
  TXSEQUENCE0,
  TXSEQUENCE1,
  TXSEQUENCE2,
  TXSEQUENCE3,
  TXSEQUENCE4,
  TXSEQUENCE5,
  TXSEQUENCE6,
  TXSEQUENCE7,
  TXSLEWCTRL0,
  TXSLEWCTRL1,
  TXSLEWCTRL2,
  TXSLEWCTRL3,
  TXSLEWCTRL4,
  TXSLEWCTRL5,
  TXSLEWCTRL6,
  TXSLEWCTRL7,
  TXUSRCLK0,
  TXUSRCLK1,
  TXUSRCLK2,
  TXUSRCLK3,
  TXUSRCLK4,
  TXUSRCLK5,
  TXUSRCLK6,
  TXUSRCLK7
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CFGCLK ;
input CFGDATAVALID ;
input CFGREADBACKB ;
input DRPCLK0 ;
input DRPCLK1 ;
input DRPCLKSEL ;
input DRPEN ;
input DRPWE ;
input FARLOOPBACKEN0 ;
input FARLOOPBACKEN1 ;
input FARLOOPBACKEN2 ;
input FARLOOPBACKEN3 ;
input FARLOOPBACKEN4 ;
input FARLOOPBACKEN5 ;
input FARLOOPBACKEN6 ;
input FARLOOPBACKEN7 ;
input GTREFCLK0N ;
input GTREFCLK0P ;
input GTREFCLK1N ;
input GTREFCLK1P ;
input GTZINIT ;
input GTZRXN0 ;
input GTZRXN1 ;
input GTZRXN2 ;
input GTZRXN3 ;
input GTZRXN4 ;
input GTZRXN5 ;
input GTZRXN6 ;
input GTZRXN7 ;
input GTZRXP0 ;
input GTZRXP1 ;
input GTZRXP2 ;
input GTZRXP3 ;
input GTZRXP4 ;
input GTZRXP5 ;
input GTZRXP6 ;
input GTZRXP7 ;
input GTZRXRESET0 ;
input GTZRXRESET1 ;
input GTZRXRESET2 ;
input GTZRXRESET3 ;
input GTZRXRESET4 ;
input GTZRXRESET5 ;
input GTZRXRESET6 ;
input GTZRXRESET7 ;
input GTZTXRESET0 ;
input GTZTXRESET1 ;
input GTZTXRESET2 ;
input GTZTXRESET3 ;
input GTZTXRESET4 ;
input GTZTXRESET5 ;
input GTZTXRESET6 ;
input GTZTXRESET7 ;
input NEARLOOPBACKEN0 ;
input NEARLOOPBACKEN1 ;
input NEARLOOPBACKEN2 ;
input NEARLOOPBACKEN3 ;
input NEARLOOPBACKEN4 ;
input NEARLOOPBACKEN5 ;
input NEARLOOPBACKEN6 ;
input NEARLOOPBACKEN7 ;
input PLLRECALEN0 ;
input PLLRECALEN1 ;
input PLLRECALEN2 ;
input PLLRECALEN3 ;
input PLLRECALEN4 ;
input PLLRECALEN5 ;
input PLLRECALEN6 ;
input PLLRECALEN7 ;
input REFCLKSEL0 ;
input REFCLKSEL1 ;
input REFCLKSEL2 ;
input REFCLKSEL3 ;
input REFCLKSEL4 ;
input REFCLKSEL5 ;
input REFCLKSEL6 ;
input REFCLKSEL7 ;
input RXBITSLIP0 ;
input RXBITSLIP1 ;
input RXBITSLIP2 ;
input RXBITSLIP3 ;
input RXBITSLIP4 ;
input RXBITSLIP5 ;
input RXBITSLIP6 ;
input RXBITSLIP7 ;
input RXEN0 ;
input RXEN1 ;
input RXEN2 ;
input RXEN3 ;
input RXEN4 ;
input RXEN5 ;
input RXEN6 ;
input RXEN7 ;
input RXFIBRESET0 ;
input RXFIBRESET1 ;
input RXFIBRESET2 ;
input RXFIBRESET3 ;
input RXFIBRESET4 ;
input RXFIBRESET5 ;
input RXFIBRESET6 ;
input RXFIBRESET7 ;
input RXLATCLK ;
input RXPOLARITY0 ;
input RXPOLARITY1 ;
input RXPOLARITY2 ;
input RXPOLARITY3 ;
input RXPOLARITY4 ;
input RXPOLARITY5 ;
input RXPOLARITY6 ;
input RXPOLARITY7 ;
input RXPRBSEN0 ;
input RXPRBSEN1 ;
input RXPRBSEN2 ;
input RXPRBSEN3 ;
input RXPRBSEN4 ;
input RXPRBSEN5 ;
input RXPRBSEN6 ;
input RXPRBSEN7 ;
input RXUSRCLK0 ;
input RXUSRCLK1 ;
input RXUSRCLK2 ;
input RXUSRCLK3 ;
input RXUSRCLK4 ;
input RXUSRCLK5 ;
input RXUSRCLK6 ;
input RXUSRCLK7 ;
input SBUSCLKSEL ;
input SBUSRESETB ;
input SPARESBUSEXECUTEB ;
input SPARESBUSRCVDATAVALIDSEL ;
input TSTRSVD0 ;
input TSTRSVD1 ;
input TSTRSVD2 ;
input TSTRSVD3 ;
input TXEN0 ;
input TXEN1 ;
input TXEN2 ;
input TXEN3 ;
input TXEN4 ;
input TXEN5 ;
input TXEN6 ;
input TXEN7 ;
input TXFIBRESET0 ;
input TXFIBRESET1 ;
input TXFIBRESET2 ;
input TXFIBRESET3 ;
input TXFIBRESET4 ;
input TXFIBRESET5 ;
input TXFIBRESET6 ;
input TXFIBRESET7 ;
input TXLATCLK ;
input TXOUTPUTEN0 ;
input TXOUTPUTEN1 ;
input TXOUTPUTEN2 ;
input TXOUTPUTEN3 ;
input TXOUTPUTEN4 ;
input TXOUTPUTEN5 ;
input TXOUTPUTEN6 ;
input TXOUTPUTEN7 ;
input TXOVERRIDEEN0 ;
input TXOVERRIDEEN1 ;
input TXOVERRIDEEN2 ;
input TXOVERRIDEEN3 ;
input TXOVERRIDEEN4 ;
input TXOVERRIDEEN5 ;
input TXOVERRIDEEN6 ;
input TXOVERRIDEEN7 ;
input TXOVERRIDEIN0 ;
input TXOVERRIDEIN1 ;
input TXOVERRIDEIN2 ;
input TXOVERRIDEIN3 ;
input TXOVERRIDEIN4 ;
input TXOVERRIDEIN5 ;
input TXOVERRIDEIN6 ;
input TXOVERRIDEIN7 ;
input TXPHASECALEN0 ;
input TXPHASECALEN1 ;
input TXPHASECALEN2 ;
input TXPHASECALEN3 ;
input TXPHASECALEN4 ;
input TXPHASECALEN5 ;
input TXPHASECALEN6 ;
input TXPHASECALEN7 ;
input TXPHASESLIP0 ;
input TXPHASESLIP1 ;
input TXPHASESLIP2 ;
input TXPHASESLIP3 ;
input TXPHASESLIP4 ;
input TXPHASESLIP5 ;
input TXPHASESLIP6 ;
input TXPHASESLIP7 ;
input TXPOLARITY0 ;
input TXPOLARITY1 ;
input TXPOLARITY2 ;
input TXPOLARITY3 ;
input TXPOLARITY4 ;
input TXPOLARITY5 ;
input TXPOLARITY6 ;
input TXPOLARITY7 ;
input TXPRBSEN0 ;
input TXPRBSEN1 ;
input TXPRBSEN2 ;
input TXPRBSEN3 ;
input TXPRBSEN4 ;
input TXPRBSEN5 ;
input TXPRBSEN6 ;
input TXPRBSEN7 ;
input TXUSRCLK0 ;
input TXUSRCLK1 ;
input TXUSRCLK2 ;
input TXUSRCLK3 ;
input TXUSRCLK4 ;
input TXUSRCLK5 ;
input TXUSRCLK6 ;
input TXUSRCLK7 ;
input [14:0] RSVDIN ;
input [159:0] TXDATA0 ;
input [159:0] TXDATA1 ;
input [159:0] TXDATA2 ;
input [159:0] TXDATA3 ;
input [159:0] TXDATA4 ;
input [159:0] TXDATA5 ;
input [159:0] TXDATA6 ;
input [159:0] TXDATA7 ;
input [15:0] CORECNTL0 ;
input [15:0] CORECNTL1 ;
input [15:0] CORECNTL2 ;
input [15:0] CORECNTL3 ;
input [15:0] CORECNTL4 ;
input [15:0] CORECNTL5 ;
input [15:0] CORECNTL6 ;
input [15:0] CORECNTL7 ;
input [15:0] DRPADDR ;
input [1:0] CFGFORCESEUERRB ;
input [1:0] RXDATAWIDTH0 ;
input [1:0] RXDATAWIDTH1 ;
input [1:0] RXDATAWIDTH2 ;
input [1:0] RXDATAWIDTH3 ;
input [1:0] RXDATAWIDTH4 ;
input [1:0] RXDATAWIDTH5 ;
input [1:0] RXDATAWIDTH6 ;
input [1:0] RXDATAWIDTH7 ;
input [1:0] TXDATAWIDTH0 ;
input [1:0] TXDATAWIDTH1 ;
input [1:0] TXDATAWIDTH2 ;
input [1:0] TXDATAWIDTH3 ;
input [1:0] TXDATAWIDTH4 ;
input [1:0] TXDATAWIDTH5 ;
input [1:0] TXDATAWIDTH6 ;
input [1:0] TXDATAWIDTH7 ;
input [1:0] TXSLEWCTRL0 ;
input [1:0] TXSLEWCTRL1 ;
input [1:0] TXSLEWCTRL2 ;
input [1:0] TXSLEWCTRL3 ;
input [1:0] TXSLEWCTRL4 ;
input [1:0] TXSLEWCTRL5 ;
input [1:0] TXSLEWCTRL6 ;
input [1:0] TXSLEWCTRL7 ;
input [2:0] CFGDEBUGMODEB ;
input [2:0] FIBRSVDIN0 ;
input [2:0] FIBRSVDIN1 ;
input [2:0] FIBRSVDIN2 ;
input [2:0] FIBRSVDIN3 ;
input [2:0] FIBRSVDIN4 ;
input [2:0] FIBRSVDIN5 ;
input [2:0] FIBRSVDIN6 ;
input [2:0] FIBRSVDIN7 ;
input [2:0] RXPRBSSEL0 ;
input [2:0] RXPRBSSEL1 ;
input [2:0] RXPRBSSEL2 ;
input [2:0] RXPRBSSEL3 ;
input [2:0] RXPRBSSEL4 ;
input [2:0] RXPRBSSEL5 ;
input [2:0] RXPRBSSEL6 ;
input [2:0] RXPRBSSEL7 ;
input [2:0] TXPRBSSEL0 ;
input [2:0] TXPRBSSEL1 ;
input [2:0] TXPRBSSEL2 ;
input [2:0] TXPRBSSEL3 ;
input [2:0] TXPRBSSEL4 ;
input [2:0] TXPRBSSEL5 ;
input [2:0] TXPRBSSEL6 ;
input [2:0] TXPRBSSEL7 ;
input [31:0] CFGDATA ;
input [31:0] DRPDI ;
input [31:0] SPARESBUSDATA ;
input [3:0] TXEQPRECTRL0 ;
input [3:0] TXEQPRECTRL1 ;
input [3:0] TXEQPRECTRL2 ;
input [3:0] TXEQPRECTRL3 ;
input [3:0] TXEQPRECTRL4 ;
input [3:0] TXEQPRECTRL5 ;
input [3:0] TXEQPRECTRL6 ;
input [3:0] TXEQPRECTRL7 ;
input [4:0] RXGEARBOXSLIP0 ;
input [4:0] RXGEARBOXSLIP1 ;
input [4:0] RXGEARBOXSLIP2 ;
input [4:0] RXGEARBOXSLIP3 ;
input [4:0] RXGEARBOXSLIP4 ;
input [4:0] RXGEARBOXSLIP5 ;
input [4:0] RXGEARBOXSLIP6 ;
input [4:0] RXGEARBOXSLIP7 ;
input [6:0] TXSEQUENCE0 ;
input [6:0] TXSEQUENCE1 ;
input [6:0] TXSEQUENCE2 ;
input [6:0] TXSEQUENCE3 ;
input [6:0] TXSEQUENCE4 ;
input [6:0] TXSEQUENCE5 ;
input [6:0] TXSEQUENCE6 ;
input [6:0] TXSEQUENCE7 ;
input [7:0] REFSEL0 ;
input [7:0] REFSEL1 ;
input [7:0] REFSEL2 ;
input [7:0] REFSEL3 ;
input [7:0] REFSEL4 ;
input [7:0] REFSEL5 ;
input [7:0] REFSEL6 ;
input [7:0] REFSEL7 ;
input [7:0] SPARESBUSCOMMAND ;
input [7:0] SPARESBUSDATAADDR ;
input [7:0] SPARESBUSRECADDR ;
input [7:0] TXATTNCTRL0 ;
input [7:0] TXATTNCTRL1 ;
input [7:0] TXATTNCTRL2 ;
input [7:0] TXATTNCTRL3 ;
input [7:0] TXATTNCTRL4 ;
input [7:0] TXATTNCTRL5 ;
input [7:0] TXATTNCTRL6 ;
input [7:0] TXATTNCTRL7 ;
input [7:0] TXEQPOSTCTRL0 ;
input [7:0] TXEQPOSTCTRL1 ;
input [7:0] TXEQPOSTCTRL2 ;
input [7:0] TXEQPOSTCTRL3 ;
input [7:0] TXEQPOSTCTRL4 ;
input [7:0] TXEQPOSTCTRL5 ;
input [7:0] TXEQPOSTCTRL6 ;
input [7:0] TXEQPOSTCTRL7 ;
input [8:0] RXRATESEL0 ;
input [8:0] RXRATESEL1 ;
input [8:0] RXRATESEL2 ;
input [8:0] RXRATESEL3 ;
input [8:0] RXRATESEL4 ;
input [8:0] RXRATESEL5 ;
input [8:0] RXRATESEL6 ;
input [8:0] RXRATESEL7 ;
input [8:0] TXRATESEL0 ;
input [8:0] TXRATESEL1 ;
input [8:0] TXRATESEL2 ;
input [8:0] TXRATESEL3 ;
input [8:0] TXRATESEL4 ;
input [8:0] TXRATESEL5 ;
input [8:0] TXRATESEL6 ;
input [8:0] TXRATESEL7 ;
input [9:0] TSTRSVD4 ;
input [9:0] TXHEADER0 ;
input [9:0] TXHEADER1 ;
input [9:0] TXHEADER2 ;
input [9:0] TXHEADER3 ;
input [9:0] TXHEADER4 ;
input [9:0] TXHEADER5 ;
input [9:0] TXHEADER6 ;
input [9:0] TXHEADER7 ;
output CFGBADVERSIONB ;
output CFGGTZDONEB ;
output DRPRDY ;
output DRPWDTERR ;
output GTZINITDONEB ;
output GTZTXN0 ;
output GTZTXN1 ;
output GTZTXN2 ;
output GTZTXN3 ;
output GTZTXN4 ;
output GTZTXN5 ;
output GTZTXN6 ;
output GTZTXN7 ;
output GTZTXP0 ;
output GTZTXP1 ;
output GTZTXP2 ;
output GTZTXP3 ;
output GTZTXP4 ;
output GTZTXP5 ;
output GTZTXP6 ;
output GTZTXP7 ;
output RXOUTCLK0 ;
output RXOUTCLK1 ;
output RXOUTCLK2 ;
output RXOUTCLK3 ;
output RXPRBSPASS0 ;
output RXPRBSPASS1 ;
output RXPRBSPASS2 ;
output RXPRBSPASS3 ;
output RXPRBSPASS4 ;
output RXPRBSPASS5 ;
output RXPRBSPASS6 ;
output RXPRBSPASS7 ;
output RXRDY0 ;
output RXRDY1 ;
output RXRDY2 ;
output RXRDY3 ;
output RXRDY4 ;
output RXRDY5 ;
output RXRDY6 ;
output RXRDY7 ;
output RXRESETDONE0 ;
output RXRESETDONE1 ;
output RXRESETDONE2 ;
output RXRESETDONE3 ;
output RXRESETDONE4 ;
output RXRESETDONE5 ;
output RXRESETDONE6 ;
output RXRESETDONE7 ;
output RXSIGNALOK0 ;
output RXSIGNALOK1 ;
output RXSIGNALOK2 ;
output RXSIGNALOK3 ;
output RXSIGNALOK4 ;
output RXSIGNALOK5 ;
output RXSIGNALOK6 ;
output RXSIGNALOK7 ;
output SPARESBUSDONE ;
output SPARESBUSRCVDATAVALID ;
output TXOUTCLK0 ;
output TXOUTCLK1 ;
output TXRDY0 ;
output TXRDY1 ;
output TXRDY2 ;
output TXRDY3 ;
output TXRDY4 ;
output TXRDY5 ;
output TXRDY6 ;
output TXRDY7 ;
output TXRESETDONE0 ;
output TXRESETDONE1 ;
output TXRESETDONE2 ;
output TXRESETDONE3 ;
output TXRESETDONE4 ;
output TXRESETDONE5 ;
output TXRESETDONE6 ;
output TXRESETDONE7 ;
output [159:0] RXDATA0 ;
output [159:0] RXDATA1 ;
output [159:0] RXDATA2 ;
output [159:0] RXDATA3 ;
output [159:0] RXDATA4 ;
output [159:0] RXDATA5 ;
output [159:0] RXDATA6 ;
output [159:0] RXDATA7 ;
output [15:0] RSVDOUT ;
output [1:0] CFGCRCERRB ;
output [1:0] CFGSEUERRB ;
output [1:0] RXFIFOSTATUS0 ;
output [1:0] RXFIFOSTATUS1 ;
output [1:0] RXFIFOSTATUS2 ;
output [1:0] RXFIFOSTATUS3 ;
output [1:0] RXFIFOSTATUS4 ;
output [1:0] RXFIFOSTATUS5 ;
output [1:0] RXFIFOSTATUS6 ;
output [1:0] RXFIFOSTATUS7 ;
output [1:0] TXFIFOSTATUS0 ;
output [1:0] TXFIFOSTATUS1 ;
output [1:0] TXFIFOSTATUS2 ;
output [1:0] TXFIFOSTATUS3 ;
output [1:0] TXFIFOSTATUS4 ;
output [1:0] TXFIFOSTATUS5 ;
output [1:0] TXFIFOSTATUS6 ;
output [1:0] TXFIFOSTATUS7 ;
output [2:0] DRPSTATUS ;
output [2:0] SPARESBUSRESULTCODE ;
output [31:0] DRPDO ;
output [31:0] SPARESBUSDATAOUT ;
output [3:0] FIBRSVDOUT0 ;
output [3:0] FIBRSVDOUT1 ;
output [3:0] FIBRSVDOUT2 ;
output [3:0] FIBRSVDOUT3 ;
output [3:0] FIBRSVDOUT4 ;
output [3:0] FIBRSVDOUT5 ;
output [3:0] FIBRSVDOUT6 ;
output [3:0] FIBRSVDOUT7 ;
output [4:0] RXDATAVALID0 ;
output [4:0] RXDATAVALID1 ;
output [4:0] RXDATAVALID2 ;
output [4:0] RXDATAVALID3 ;
output [4:0] RXDATAVALID4 ;
output [4:0] RXDATAVALID5 ;
output [4:0] RXDATAVALID6 ;
output [4:0] RXDATAVALID7 ;
output [4:0] RXHEADERVALID0 ;
output [4:0] RXHEADERVALID1 ;
output [4:0] RXHEADERVALID2 ;
output [4:0] RXHEADERVALID3 ;
output [4:0] RXHEADERVALID4 ;
output [4:0] RXHEADERVALID5 ;
output [4:0] RXHEADERVALID6 ;
output [4:0] RXHEADERVALID7 ;
output [4:0] TXPHASEOUT0 ;
output [4:0] TXPHASEOUT1 ;
output [4:0] TXPHASEOUT2 ;
output [4:0] TXPHASEOUT3 ;
output [4:0] TXPHASEOUT4 ;
output [4:0] TXPHASEOUT5 ;
output [4:0] TXPHASEOUT6 ;
output [4:0] TXPHASEOUT7 ;
output [9:0] RXHEADER0 ;
output [9:0] RXHEADER1 ;
output [9:0] RXHEADER2 ;
output [9:0] RXHEADER3 ;
output [9:0] RXHEADER4 ;
output [9:0] RXHEADER5 ;
output [9:0] RXHEADER6 ;
output [9:0] RXHEADER7 ;
parameter [0:0] ACCLK_HYST_EN_0 = 1'b0;
parameter [0:0] ACCLK_HYST_EN_1 = 1'b0;
parameter [0:0] ACCLK_MUX_DIV2_SEL_0 = 1'b1;
parameter [0:0] ACCLK_MUX_DIV2_SEL_1 = 1'b1;
parameter [0:0] ACCLK_TERM_EN_0 = 1'b0;
parameter [0:0] ACCLK_TERM_EN_1 = 1'b0;
parameter [31:0] BROADCAST_CTRL_LANE0 = 32'h00000000;
parameter [31:0] BROADCAST_CTRL_LANE1 = 32'h00000000;
parameter [31:0] BROADCAST_CTRL_LANE2 = 32'h00000000;
parameter [31:0] BROADCAST_CTRL_LANE3 = 32'h00000000;
parameter [31:0] BROADCAST_CTRL_LANE4 = 32'h00000000;
parameter [31:0] BROADCAST_CTRL_LANE5 = 32'h00000000;
parameter [31:0] BROADCAST_CTRL_LANE6 = 32'h00000000;
parameter [31:0] BROADCAST_CTRL_LANE7 = 32'h00000000;
parameter [0:0] BYPASS_FIRMWARE_CRC_CHECK = 1'b0;
parameter [1:0] BYPASS_SERDES_CONFIG = 2'b00;
parameter [0:0] CONFIG_MEM_WRITE_EN = 1'b0;
parameter [1:0] DRV_IMP_CONFIG_LANE0 = 2'b01;
parameter [1:0] DRV_IMP_CONFIG_LANE1 = 2'b01;
parameter [1:0] DRV_IMP_CONFIG_LANE2 = 2'b01;
parameter [1:0] DRV_IMP_CONFIG_LANE3 = 2'b01;
parameter [1:0] DRV_IMP_CONFIG_LANE4 = 2'b01;
parameter [1:0] DRV_IMP_CONFIG_LANE5 = 2'b01;
parameter [1:0] DRV_IMP_CONFIG_LANE6 = 2'b01;
parameter [1:0] DRV_IMP_CONFIG_LANE7 = 2'b01;
parameter [16:0] FIB_ASYNC_CTRL_LANE0 = 17'h0FDFF;
parameter [16:0] FIB_ASYNC_CTRL_LANE1 = 17'h0FDFF;
parameter [16:0] FIB_ASYNC_CTRL_LANE2 = 17'h0FDFF;
parameter [16:0] FIB_ASYNC_CTRL_LANE3 = 17'h0FDFF;
parameter [16:0] FIB_ASYNC_CTRL_LANE4 = 17'h0FDFF;
parameter [16:0] FIB_ASYNC_CTRL_LANE5 = 17'h0FDFF;
parameter [16:0] FIB_ASYNC_CTRL_LANE6 = 17'h0FDFF;
parameter [16:0] FIB_ASYNC_CTRL_LANE7 = 17'h0FDFF;
parameter FIB_IGNORE_BROADCAST_LANE0 = "FALSE";
parameter FIB_IGNORE_BROADCAST_LANE1 = "FALSE";
parameter FIB_IGNORE_BROADCAST_LANE2 = "FALSE";
parameter FIB_IGNORE_BROADCAST_LANE3 = "FALSE";
parameter FIB_IGNORE_BROADCAST_LANE4 = "FALSE";
parameter FIB_IGNORE_BROADCAST_LANE5 = "FALSE";
parameter FIB_IGNORE_BROADCAST_LANE6 = "FALSE";
parameter FIB_IGNORE_BROADCAST_LANE7 = "FALSE";
parameter FIB_LOOPBACK_SEL_LANE0 = "NORMAL";
parameter FIB_LOOPBACK_SEL_LANE1 = "NORMAL";
parameter FIB_LOOPBACK_SEL_LANE2 = "NORMAL";
parameter FIB_LOOPBACK_SEL_LANE3 = "NORMAL";
parameter FIB_LOOPBACK_SEL_LANE4 = "NORMAL";
parameter FIB_LOOPBACK_SEL_LANE5 = "NORMAL";
parameter FIB_LOOPBACK_SEL_LANE6 = "NORMAL";
parameter FIB_LOOPBACK_SEL_LANE7 = "NORMAL";
parameter [7:0] FIB_MULTICAST_GROUP_ID_LANE0 = 8'h00;
parameter [7:0] FIB_MULTICAST_GROUP_ID_LANE1 = 8'h00;
parameter [7:0] FIB_MULTICAST_GROUP_ID_LANE2 = 8'h00;
parameter [7:0] FIB_MULTICAST_GROUP_ID_LANE3 = 8'h00;
parameter [7:0] FIB_MULTICAST_GROUP_ID_LANE4 = 8'h00;
parameter [7:0] FIB_MULTICAST_GROUP_ID_LANE5 = 8'h00;
parameter [7:0] FIB_MULTICAST_GROUP_ID_LANE6 = 8'h00;
parameter [7:0] FIB_MULTICAST_GROUP_ID_LANE7 = 8'h00;
parameter FIB_NEAREND_LPBK_CLK_SEL_LANE0 = "TXOUTCLKPMA";
parameter FIB_NEAREND_LPBK_CLK_SEL_LANE1 = "TXOUTCLKPMA";
parameter FIB_NEAREND_LPBK_CLK_SEL_LANE2 = "TXOUTCLKPMA";
parameter FIB_NEAREND_LPBK_CLK_SEL_LANE3 = "TXOUTCLKPMA";
parameter FIB_NEAREND_LPBK_CLK_SEL_LANE4 = "TXOUTCLKPMA";
parameter FIB_NEAREND_LPBK_CLK_SEL_LANE5 = "TXOUTCLKPMA";
parameter FIB_NEAREND_LPBK_CLK_SEL_LANE6 = "TXOUTCLKPMA";
parameter FIB_NEAREND_LPBK_CLK_SEL_LANE7 = "TXOUTCLKPMA";
parameter [31:0] FIB_RSVD_REG_LANE0 = 32'h00000000;
parameter [31:0] FIB_RSVD_REG_LANE1 = 32'h00000000;
parameter [31:0] FIB_RSVD_REG_LANE2 = 32'h00000000;
parameter [31:0] FIB_RSVD_REG_LANE3 = 32'h00000000;
parameter [31:0] FIB_RSVD_REG_LANE4 = 32'h00000000;
parameter [31:0] FIB_RSVD_REG_LANE5 = 32'h00000000;
parameter [31:0] FIB_RSVD_REG_LANE6 = 32'h00000000;
parameter [31:0] FIB_RSVD_REG_LANE7 = 32'h00000000;
parameter [0:0] GTZ_POWER_UP_LANE0 = 1'b1;
parameter [0:0] GTZ_POWER_UP_LANE1 = 1'b1;
parameter [0:0] GTZ_POWER_UP_LANE2 = 1'b1;
parameter [0:0] GTZ_POWER_UP_LANE3 = 1'b1;
parameter [0:0] GTZ_POWER_UP_LANE4 = 1'b1;
parameter [0:0] GTZ_POWER_UP_LANE5 = 1'b1;
parameter [0:0] GTZ_POWER_UP_LANE6 = 1'b1;
parameter [0:0] GTZ_POWER_UP_LANE7 = 1'b1;
parameter [0:0] IGNORE_DOUBLE_SEU_ERR = 1'b0;
parameter [0:0] IGNORE_FIRMWARE_CRC = 1'b0;
parameter [0:0] IGNORE_SINGLE_SEU_ERR = 1'b0;
parameter [4:0] MULTI_LANE_MODE = 5'b10011;
parameter [31:0] PMA_CTRL_1_LANE0 = 32'h00000000;
parameter [31:0] PMA_CTRL_1_LANE1 = 32'h00000000;
parameter [31:0] PMA_CTRL_1_LANE2 = 32'h00000000;
parameter [31:0] PMA_CTRL_1_LANE3 = 32'h00000000;
parameter [31:0] PMA_CTRL_1_LANE4 = 32'h00000000;
parameter [31:0] PMA_CTRL_1_LANE5 = 32'h00000000;
parameter [31:0] PMA_CTRL_1_LANE6 = 32'h00000000;
parameter [31:0] PMA_CTRL_1_LANE7 = 32'h00000000;
parameter [31:0] PMA_CTRL_2_LANE0 = 32'h00000000;
parameter [31:0] PMA_CTRL_2_LANE1 = 32'h00000000;
parameter [31:0] PMA_CTRL_2_LANE2 = 32'h00000000;
parameter [31:0] PMA_CTRL_2_LANE3 = 32'h00000000;
parameter [31:0] PMA_CTRL_2_LANE4 = 32'h00000000;
parameter [31:0] PMA_CTRL_2_LANE5 = 32'h00000000;
parameter [31:0] PMA_CTRL_2_LANE6 = 32'h00000000;
parameter [31:0] PMA_CTRL_2_LANE7 = 32'h00000000;
parameter [31:0] PMA_WIDTH_CTRL_LANE0 = 32'h00000000;
parameter [31:0] PMA_WIDTH_CTRL_LANE1 = 32'h00000000;
parameter [31:0] PMA_WIDTH_CTRL_LANE2 = 32'h00000000;
parameter [31:0] PMA_WIDTH_CTRL_LANE3 = 32'h00000000;
parameter [31:0] PMA_WIDTH_CTRL_LANE4 = 32'h00000000;
parameter [31:0] PMA_WIDTH_CTRL_LANE5 = 32'h00000000;
parameter [31:0] PMA_WIDTH_CTRL_LANE6 = 32'h00000000;
parameter [31:0] PMA_WIDTH_CTRL_LANE7 = 32'h00000000;
parameter [1:0] RESETDONE_IGNORE_RDY_LANE0 = 2'b00;
parameter [1:0] RESETDONE_IGNORE_RDY_LANE1 = 2'b00;
parameter [1:0] RESETDONE_IGNORE_RDY_LANE2 = 2'b00;
parameter [1:0] RESETDONE_IGNORE_RDY_LANE3 = 2'b00;
parameter [1:0] RESETDONE_IGNORE_RDY_LANE4 = 2'b00;
parameter [1:0] RESETDONE_IGNORE_RDY_LANE5 = 2'b00;
parameter [1:0] RESETDONE_IGNORE_RDY_LANE6 = 2'b00;
parameter [1:0] RESETDONE_IGNORE_RDY_LANE7 = 2'b00;
parameter [1:0] RESET_IGNORE_FIBINITDONE_LANE0 = 2'b00;
parameter [1:0] RESET_IGNORE_FIBINITDONE_LANE1 = 2'b00;
parameter [1:0] RESET_IGNORE_FIBINITDONE_LANE2 = 2'b00;
parameter [1:0] RESET_IGNORE_FIBINITDONE_LANE3 = 2'b00;
parameter [1:0] RESET_IGNORE_FIBINITDONE_LANE4 = 2'b00;
parameter [1:0] RESET_IGNORE_FIBINITDONE_LANE5 = 2'b00;
parameter [1:0] RESET_IGNORE_FIBINITDONE_LANE6 = 2'b00;
parameter [1:0] RESET_IGNORE_FIBINITDONE_LANE7 = 2'b00;
parameter [1:0] RESET_IGNORE_GTZINITDONE_LANE0 = 2'b00;
parameter [1:0] RESET_IGNORE_GTZINITDONE_LANE1 = 2'b00;
parameter [1:0] RESET_IGNORE_GTZINITDONE_LANE2 = 2'b00;
parameter [1:0] RESET_IGNORE_GTZINITDONE_LANE3 = 2'b00;
parameter [1:0] RESET_IGNORE_GTZINITDONE_LANE4 = 2'b00;
parameter [1:0] RESET_IGNORE_GTZINITDONE_LANE5 = 2'b00;
parameter [1:0] RESET_IGNORE_GTZINITDONE_LANE6 = 2'b00;
parameter [1:0] RESET_IGNORE_GTZINITDONE_LANE7 = 2'b00;
parameter [1:0] RESET_MODE_LANE0 = 2'b00;
parameter [1:0] RESET_MODE_LANE1 = 2'b00;
parameter [1:0] RESET_MODE_LANE2 = 2'b00;
parameter [1:0] RESET_MODE_LANE3 = 2'b00;
parameter [1:0] RESET_MODE_LANE4 = 2'b00;
parameter [1:0] RESET_MODE_LANE5 = 2'b00;
parameter [1:0] RESET_MODE_LANE6 = 2'b00;
parameter [1:0] RESET_MODE_LANE7 = 2'b00;
parameter [31:0] RSVD_REG_1 = 32'h00000001;
parameter [31:0] RSVD_REG_2 = 32'h00000000;
parameter [5:0] RXFIFO_BITSLIP_RESET_TIME_LANE0 = 6'h16;
parameter [5:0] RXFIFO_BITSLIP_RESET_TIME_LANE1 = 6'h16;
parameter [5:0] RXFIFO_BITSLIP_RESET_TIME_LANE2 = 6'h16;
parameter [5:0] RXFIFO_BITSLIP_RESET_TIME_LANE3 = 6'h16;
parameter [5:0] RXFIFO_BITSLIP_RESET_TIME_LANE4 = 6'h16;
parameter [5:0] RXFIFO_BITSLIP_RESET_TIME_LANE5 = 6'h16;
parameter [5:0] RXFIFO_BITSLIP_RESET_TIME_LANE6 = 6'h16;
parameter [5:0] RXFIFO_BITSLIP_RESET_TIME_LANE7 = 6'h16;
parameter RXFIFO_EN_LANE0 = "TRUE";
parameter RXFIFO_EN_LANE1 = "TRUE";
parameter RXFIFO_EN_LANE2 = "TRUE";
parameter RXFIFO_EN_LANE3 = "TRUE";
parameter RXFIFO_EN_LANE4 = "TRUE";
parameter RXFIFO_EN_LANE5 = "TRUE";
parameter RXFIFO_EN_LANE6 = "TRUE";
parameter RXFIFO_EN_LANE7 = "TRUE";
parameter RXFIFO_RESET_ON_BITSLIP_LANE0 = "TRUE";
parameter RXFIFO_RESET_ON_BITSLIP_LANE1 = "TRUE";
parameter RXFIFO_RESET_ON_BITSLIP_LANE2 = "TRUE";
parameter RXFIFO_RESET_ON_BITSLIP_LANE3 = "TRUE";
parameter RXFIFO_RESET_ON_BITSLIP_LANE4 = "TRUE";
parameter RXFIFO_RESET_ON_BITSLIP_LANE5 = "TRUE";
parameter RXFIFO_RESET_ON_BITSLIP_LANE6 = "TRUE";
parameter RXFIFO_RESET_ON_BITSLIP_LANE7 = "TRUE";
parameter RXOUTCLK0_LANE_SEL = "LANE0";
parameter RXOUTCLK1_LANE_SEL = "LANE0";
parameter RXOUTCLK2_LANE_SEL = "LANE0";
parameter RXOUTCLK3_LANE_SEL = "LANE0";
parameter RXOUTCLK_SEL_LANE0 = "RXRECCLKPMA_DIV4";
parameter RXOUTCLK_SEL_LANE1 = "RXRECCLKPMA_DIV4";
parameter RXOUTCLK_SEL_LANE2 = "RXRECCLKPMA_DIV4";
parameter RXOUTCLK_SEL_LANE3 = "RXRECCLKPMA_DIV4";
parameter RXOUTCLK_SEL_LANE4 = "RXRECCLKPMA_DIV4";
parameter RXOUTCLK_SEL_LANE5 = "RXRECCLKPMA_DIV4";
parameter RXOUTCLK_SEL_LANE6 = "RXRECCLKPMA_DIV4";
parameter RXOUTCLK_SEL_LANE7 = "RXRECCLKPMA_DIV4";
parameter [7:0] RXPMARESET_TIME_LANE0 = 8'h32;
parameter [7:0] RXPMARESET_TIME_LANE1 = 8'h32;
parameter [7:0] RXPMARESET_TIME_LANE2 = 8'h32;
parameter [7:0] RXPMARESET_TIME_LANE3 = 8'h32;
parameter [7:0] RXPMARESET_TIME_LANE4 = 8'h32;
parameter [7:0] RXPMARESET_TIME_LANE5 = 8'h32;
parameter [7:0] RXPMARESET_TIME_LANE6 = 8'h32;
parameter [7:0] RXPMARESET_TIME_LANE7 = 8'h32;
parameter [10:0] RXRESETDONE_TIME_LANE0 = 11'h21A;
parameter [10:0] RXRESETDONE_TIME_LANE1 = 11'h21A;
parameter [10:0] RXRESETDONE_TIME_LANE2 = 11'h21A;
parameter [10:0] RXRESETDONE_TIME_LANE3 = 11'h21A;
parameter [10:0] RXRESETDONE_TIME_LANE4 = 11'h21A;
parameter [10:0] RXRESETDONE_TIME_LANE5 = 11'h21A;
parameter [10:0] RXRESETDONE_TIME_LANE6 = 11'h21A;
parameter [10:0] RXRESETDONE_TIME_LANE7 = 11'h21A;
parameter RXUSRCLK_SEL_LANE0 = "RXUSRCLK0";
parameter RXUSRCLK_SEL_LANE1 = "RXUSRCLK0";
parameter RXUSRCLK_SEL_LANE2 = "RXUSRCLK0";
parameter RXUSRCLK_SEL_LANE3 = "RXUSRCLK0";
parameter RXUSRCLK_SEL_LANE4 = "RXUSRCLK0";
parameter RXUSRCLK_SEL_LANE5 = "RXUSRCLK0";
parameter RXUSRCLK_SEL_LANE6 = "RXUSRCLK0";
parameter RXUSRCLK_SEL_LANE7 = "RXUSRCLK0";
parameter [31:0] RX_ALT_PATTERN_CTRL_LANE0 = 32'h00000000;
parameter [31:0] RX_ALT_PATTERN_CTRL_LANE1 = 32'h00000000;
parameter [31:0] RX_ALT_PATTERN_CTRL_LANE2 = 32'h00000000;
parameter [31:0] RX_ALT_PATTERN_CTRL_LANE3 = 32'h00000000;
parameter [31:0] RX_ALT_PATTERN_CTRL_LANE4 = 32'h00000000;
parameter [31:0] RX_ALT_PATTERN_CTRL_LANE5 = 32'h00000000;
parameter [31:0] RX_ALT_PATTERN_CTRL_LANE6 = 32'h00000000;
parameter [31:0] RX_ALT_PATTERN_CTRL_LANE7 = 32'h00000000;
parameter RX_CLK_GATING_EN_LANE0 = "TRUE";
parameter RX_CLK_GATING_EN_LANE1 = "TRUE";
parameter RX_CLK_GATING_EN_LANE2 = "TRUE";
parameter RX_CLK_GATING_EN_LANE3 = "TRUE";
parameter RX_CLK_GATING_EN_LANE4 = "TRUE";
parameter RX_CLK_GATING_EN_LANE5 = "TRUE";
parameter RX_CLK_GATING_EN_LANE6 = "TRUE";
parameter RX_CLK_GATING_EN_LANE7 = "TRUE";
parameter [31:0] RX_DFE_PHASE_CTRL_LANE0 = 32'h00000000;
parameter [31:0] RX_DFE_PHASE_CTRL_LANE1 = 32'h00000000;
parameter [31:0] RX_DFE_PHASE_CTRL_LANE2 = 32'h00000000;
parameter [31:0] RX_DFE_PHASE_CTRL_LANE3 = 32'h00000000;
parameter [31:0] RX_DFE_PHASE_CTRL_LANE4 = 32'h00000000;
parameter [31:0] RX_DFE_PHASE_CTRL_LANE5 = 32'h00000000;
parameter [31:0] RX_DFE_PHASE_CTRL_LANE6 = 32'h00000000;
parameter [31:0] RX_DFE_PHASE_CTRL_LANE7 = 32'h00000000;
parameter [31:0] RX_ERR_MON_CTRL_LANE0 = 32'h00000000;
parameter [31:0] RX_ERR_MON_CTRL_LANE1 = 32'h00000000;
parameter [31:0] RX_ERR_MON_CTRL_LANE2 = 32'h00000000;
parameter [31:0] RX_ERR_MON_CTRL_LANE3 = 32'h00000000;
parameter [31:0] RX_ERR_MON_CTRL_LANE4 = 32'h00000000;
parameter [31:0] RX_ERR_MON_CTRL_LANE5 = 32'h00000000;
parameter [31:0] RX_ERR_MON_CTRL_LANE6 = 32'h00000000;
parameter [31:0] RX_ERR_MON_CTRL_LANE7 = 32'h00000000;
parameter [31:0] RX_FAR_LPBK_CTRL_LANE0 = 32'h00000000;
parameter [31:0] RX_FAR_LPBK_CTRL_LANE1 = 32'h00000000;
parameter [31:0] RX_FAR_LPBK_CTRL_LANE2 = 32'h00000000;
parameter [31:0] RX_FAR_LPBK_CTRL_LANE3 = 32'h00000000;
parameter [31:0] RX_FAR_LPBK_CTRL_LANE4 = 32'h00000000;
parameter [31:0] RX_FAR_LPBK_CTRL_LANE5 = 32'h00000000;
parameter [31:0] RX_FAR_LPBK_CTRL_LANE6 = 32'h00000000;
parameter [31:0] RX_FAR_LPBK_CTRL_LANE7 = 32'h00000000;
parameter [31:0] RX_GAIN_CTRL_LANE0 = 32'h00000000;
parameter [31:0] RX_GAIN_CTRL_LANE1 = 32'h00000000;
parameter [31:0] RX_GAIN_CTRL_LANE2 = 32'h00000000;
parameter [31:0] RX_GAIN_CTRL_LANE3 = 32'h00000000;
parameter [31:0] RX_GAIN_CTRL_LANE4 = 32'h00000000;
parameter [31:0] RX_GAIN_CTRL_LANE5 = 32'h00000000;
parameter [31:0] RX_GAIN_CTRL_LANE6 = 32'h00000000;
parameter [31:0] RX_GAIN_CTRL_LANE7 = 32'h00000000;
parameter RX_MODE_SEL_LANE0 = "GB_100GBASE_R4";
parameter RX_MODE_SEL_LANE1 = "GB_100GBASE_R4";
parameter RX_MODE_SEL_LANE2 = "GB_100GBASE_R4";
parameter RX_MODE_SEL_LANE3 = "GB_100GBASE_R4";
parameter RX_MODE_SEL_LANE4 = "GB_100GBASE_R4";
parameter RX_MODE_SEL_LANE5 = "GB_100GBASE_R4";
parameter RX_MODE_SEL_LANE6 = "GB_100GBASE_R4";
parameter RX_MODE_SEL_LANE7 = "GB_100GBASE_R4";
parameter [31:0] RX_PATTERN_CTRL_LANE0 = 32'h02000000;
parameter [31:0] RX_PATTERN_CTRL_LANE1 = 32'h02000000;
parameter [31:0] RX_PATTERN_CTRL_LANE2 = 32'h02000000;
parameter [31:0] RX_PATTERN_CTRL_LANE3 = 32'h02000000;
parameter [31:0] RX_PATTERN_CTRL_LANE4 = 32'h02000000;
parameter [31:0] RX_PATTERN_CTRL_LANE5 = 32'h02000000;
parameter [31:0] RX_PATTERN_CTRL_LANE6 = 32'h02000000;
parameter [31:0] RX_PATTERN_CTRL_LANE7 = 32'h02000000;
parameter [31:0] RX_PHASE_INT_CTRL_LANE0 = 32'h00000000;
parameter [31:0] RX_PHASE_INT_CTRL_LANE1 = 32'h00000000;
parameter [31:0] RX_PHASE_INT_CTRL_LANE2 = 32'h00000000;
parameter [31:0] RX_PHASE_INT_CTRL_LANE3 = 32'h00000000;
parameter [31:0] RX_PHASE_INT_CTRL_LANE4 = 32'h00000000;
parameter [31:0] RX_PHASE_INT_CTRL_LANE5 = 32'h00000000;
parameter [31:0] RX_PHASE_INT_CTRL_LANE6 = 32'h00000000;
parameter [31:0] RX_PHASE_INT_CTRL_LANE7 = 32'h00000000;
parameter [2:0] RX_SAMPLE_PERIOD_LANE0 = 3'b110;
parameter [2:0] RX_SAMPLE_PERIOD_LANE1 = 3'b110;
parameter [2:0] RX_SAMPLE_PERIOD_LANE2 = 3'b110;
parameter [2:0] RX_SAMPLE_PERIOD_LANE3 = 3'b110;
parameter [2:0] RX_SAMPLE_PERIOD_LANE4 = 3'b110;
parameter [2:0] RX_SAMPLE_PERIOD_LANE5 = 3'b110;
parameter [2:0] RX_SAMPLE_PERIOD_LANE6 = 3'b110;
parameter [2:0] RX_SAMPLE_PERIOD_LANE7 = 3'b110;
parameter [31:0] RX_SIGNAL_OK_CTRL_LANE0 = 32'h00500000;
parameter [31:0] RX_SIGNAL_OK_CTRL_LANE1 = 32'h00500000;
parameter [31:0] RX_SIGNAL_OK_CTRL_LANE2 = 32'h00500000;
parameter [31:0] RX_SIGNAL_OK_CTRL_LANE3 = 32'h00500000;
parameter [31:0] RX_SIGNAL_OK_CTRL_LANE4 = 32'h00500000;
parameter [31:0] RX_SIGNAL_OK_CTRL_LANE5 = 32'h00500000;
parameter [31:0] RX_SIGNAL_OK_CTRL_LANE6 = 32'h00500000;
parameter [31:0] RX_SIGNAL_OK_CTRL_LANE7 = 32'h00500000;
parameter [31:0] RX_USER_REG_CTRL_LANE0 = 32'h00000000;
parameter [31:0] RX_USER_REG_CTRL_LANE1 = 32'h00000000;
parameter [31:0] RX_USER_REG_CTRL_LANE2 = 32'h00000000;
parameter [31:0] RX_USER_REG_CTRL_LANE3 = 32'h00000000;
parameter [31:0] RX_USER_REG_CTRL_LANE4 = 32'h00000000;
parameter [31:0] RX_USER_REG_CTRL_LANE5 = 32'h00000000;
parameter [31:0] RX_USER_REG_CTRL_LANE6 = 32'h00000000;
parameter [31:0] RX_USER_REG_CTRL_LANE7 = 32'h00000000;
parameter [3:0] SBUS_CLK_DIV = 4'h3;
parameter [0:0] SBUS_CLK_DIV_NON_2N_EN = 1'b0;
parameter [11:0] SBUS_CLK_DIV_NON_2N_RESET_VAL = 12'hFFF;
parameter [31:0] SBUS_OVRD_ANALOG_CTRL_LANE0 = 32'h00000000;
parameter [31:0] SBUS_OVRD_ANALOG_CTRL_LANE1 = 32'h00000000;
parameter [31:0] SBUS_OVRD_ANALOG_CTRL_LANE2 = 32'h00000000;
parameter [31:0] SBUS_OVRD_ANALOG_CTRL_LANE3 = 32'h00000000;
parameter [31:0] SBUS_OVRD_ANALOG_CTRL_LANE4 = 32'h00000000;
parameter [31:0] SBUS_OVRD_ANALOG_CTRL_LANE5 = 32'h00000000;
parameter [31:0] SBUS_OVRD_ANALOG_CTRL_LANE6 = 32'h00000000;
parameter [31:0] SBUS_OVRD_ANALOG_CTRL_LANE7 = 32'h00000000;
parameter [31:0] SBUS_OVRD_CORE_CTRL_LANE0 = 32'h00000000;
parameter [31:0] SBUS_OVRD_CORE_CTRL_LANE1 = 32'h00000000;
parameter [31:0] SBUS_OVRD_CORE_CTRL_LANE2 = 32'h00000000;
parameter [31:0] SBUS_OVRD_CORE_CTRL_LANE3 = 32'h00000000;
parameter [31:0] SBUS_OVRD_CORE_CTRL_LANE4 = 32'h00000000;
parameter [31:0] SBUS_OVRD_CORE_CTRL_LANE5 = 32'h00000000;
parameter [31:0] SBUS_OVRD_CORE_CTRL_LANE6 = 32'h00000000;
parameter [31:0] SBUS_OVRD_CORE_CTRL_LANE7 = 32'h00000000;
parameter [31:0] SBUS_TEST_RW_LANE0 = 32'h00000000;
parameter [31:0] SBUS_TEST_RW_LANE1 = 32'h00000000;
parameter [31:0] SBUS_TEST_RW_LANE2 = 32'h00000000;
parameter [31:0] SBUS_TEST_RW_LANE3 = 32'h00000000;
parameter [31:0] SBUS_TEST_RW_LANE4 = 32'h00000000;
parameter [31:0] SBUS_TEST_RW_LANE5 = 32'h00000000;
parameter [31:0] SBUS_TEST_RW_LANE6 = 32'h00000000;
parameter [31:0] SBUS_TEST_RW_LANE7 = 32'h00000000;
parameter [31:0] SERDES_CONTROL_REG_LANE0 = 32'h00000002;
parameter [31:0] SERDES_CONTROL_REG_LANE1 = 32'h00000002;
parameter [31:0] SERDES_CONTROL_REG_LANE2 = 32'h00000002;
parameter [31:0] SERDES_CONTROL_REG_LANE3 = 32'h00000002;
parameter [31:0] SERDES_CONTROL_REG_LANE4 = 32'h00000002;
parameter [31:0] SERDES_CONTROL_REG_LANE5 = 32'h00000002;
parameter [31:0] SERDES_CONTROL_REG_LANE6 = 32'h00000002;
parameter [31:0] SERDES_CONTROL_REG_LANE7 = 32'h00000002;
parameter SIM_GTZRESET_SPEEDUP = "TRUE";
parameter SIM_VERSION = "1.0";
parameter TXFIFO_EN_LANE0 = "TRUE";
parameter TXFIFO_EN_LANE1 = "TRUE";
parameter TXFIFO_EN_LANE2 = "TRUE";
parameter TXFIFO_EN_LANE3 = "TRUE";
parameter TXFIFO_EN_LANE4 = "TRUE";
parameter TXFIFO_EN_LANE5 = "TRUE";
parameter TXFIFO_EN_LANE6 = "TRUE";
parameter TXFIFO_EN_LANE7 = "TRUE";
parameter TXOUTCLK0_LANE_SEL = "LANE0";
parameter TXOUTCLK1_LANE_SEL = "LANE0";
parameter TXOUTCLK_SEL_LANE0 = "TXOUTCLKPMA_DIV4";
parameter TXOUTCLK_SEL_LANE1 = "TXOUTCLKPMA_DIV4";
parameter TXOUTCLK_SEL_LANE2 = "TXOUTCLKPMA_DIV4";
parameter TXOUTCLK_SEL_LANE3 = "TXOUTCLKPMA_DIV4";
parameter TXOUTCLK_SEL_LANE4 = "TXOUTCLKPMA_DIV4";
parameter TXOUTCLK_SEL_LANE5 = "TXOUTCLKPMA_DIV4";
parameter TXOUTCLK_SEL_LANE6 = "TXOUTCLKPMA_DIV4";
parameter TXOUTCLK_SEL_LANE7 = "TXOUTCLKPMA_DIV4";
parameter [7:0] TXPMARESET_TIME_LANE0 = 8'h32;
parameter [7:0] TXPMARESET_TIME_LANE1 = 8'h32;
parameter [7:0] TXPMARESET_TIME_LANE2 = 8'h32;
parameter [7:0] TXPMARESET_TIME_LANE3 = 8'h32;
parameter [7:0] TXPMARESET_TIME_LANE4 = 8'h32;
parameter [7:0] TXPMARESET_TIME_LANE5 = 8'h32;
parameter [7:0] TXPMARESET_TIME_LANE6 = 8'h32;
parameter [7:0] TXPMARESET_TIME_LANE7 = 8'h32;
parameter [10:0] TXRESETDONE_TIME_LANE0 = 11'h21A;
parameter [10:0] TXRESETDONE_TIME_LANE1 = 11'h21A;
parameter [10:0] TXRESETDONE_TIME_LANE2 = 11'h21A;
parameter [10:0] TXRESETDONE_TIME_LANE3 = 11'h21A;
parameter [10:0] TXRESETDONE_TIME_LANE4 = 11'h21A;
parameter [10:0] TXRESETDONE_TIME_LANE5 = 11'h21A;
parameter [10:0] TXRESETDONE_TIME_LANE6 = 11'h21A;
parameter [10:0] TXRESETDONE_TIME_LANE7 = 11'h21A;
parameter TXUSRCLK_SEL_LANE0 = "TXUSRCLK0";
parameter TXUSRCLK_SEL_LANE1 = "TXUSRCLK0";
parameter TXUSRCLK_SEL_LANE2 = "TXUSRCLK0";
parameter TXUSRCLK_SEL_LANE3 = "TXUSRCLK0";
parameter TXUSRCLK_SEL_LANE4 = "TXUSRCLK0";
parameter TXUSRCLK_SEL_LANE5 = "TXUSRCLK0";
parameter TXUSRCLK_SEL_LANE6 = "TXUSRCLK0";
parameter TXUSRCLK_SEL_LANE7 = "TXUSRCLK0";
parameter TX_CLK_GATING_EN_LANE0 = "TRUE";
parameter TX_CLK_GATING_EN_LANE1 = "TRUE";
parameter TX_CLK_GATING_EN_LANE2 = "TRUE";
parameter TX_CLK_GATING_EN_LANE3 = "TRUE";
parameter TX_CLK_GATING_EN_LANE4 = "TRUE";
parameter TX_CLK_GATING_EN_LANE5 = "TRUE";
parameter TX_CLK_GATING_EN_LANE6 = "TRUE";
parameter TX_CLK_GATING_EN_LANE7 = "TRUE";
parameter [31:0] TX_GAIN_CTRL_LANE0 = 32'h00000000;
parameter [31:0] TX_GAIN_CTRL_LANE1 = 32'h00000000;
parameter [31:0] TX_GAIN_CTRL_LANE2 = 32'h00000000;
parameter [31:0] TX_GAIN_CTRL_LANE3 = 32'h00000000;
parameter [31:0] TX_GAIN_CTRL_LANE4 = 32'h00000000;
parameter [31:0] TX_GAIN_CTRL_LANE5 = 32'h00000000;
parameter [31:0] TX_GAIN_CTRL_LANE6 = 32'h00000000;
parameter [31:0] TX_GAIN_CTRL_LANE7 = 32'h00000000;
parameter [31:0] TX_HALT_CTRL_LANE0 = 32'h00080000;
parameter [31:0] TX_HALT_CTRL_LANE1 = 32'h00080000;
parameter [31:0] TX_HALT_CTRL_LANE2 = 32'h00080000;
parameter [31:0] TX_HALT_CTRL_LANE3 = 32'h00080000;
parameter [31:0] TX_HALT_CTRL_LANE4 = 32'h00080000;
parameter [31:0] TX_HALT_CTRL_LANE5 = 32'h00080000;
parameter [31:0] TX_HALT_CTRL_LANE6 = 32'h00080000;
parameter [31:0] TX_HALT_CTRL_LANE7 = 32'h00080000;
parameter TX_MODE_SEL_LANE0 = "GB_100GBASE_R4";
parameter TX_MODE_SEL_LANE1 = "GB_100GBASE_R4";
parameter TX_MODE_SEL_LANE2 = "GB_100GBASE_R4";
parameter TX_MODE_SEL_LANE3 = "GB_100GBASE_R4";
parameter TX_MODE_SEL_LANE4 = "GB_100GBASE_R4";
parameter TX_MODE_SEL_LANE5 = "GB_100GBASE_R4";
parameter TX_MODE_SEL_LANE6 = "GB_100GBASE_R4";
parameter TX_MODE_SEL_LANE7 = "GB_100GBASE_R4";
parameter [31:0] TX_OUTPUT_CTRL_LANE0 = 32'h00000000;
parameter [31:0] TX_OUTPUT_CTRL_LANE1 = 32'h00000000;
parameter [31:0] TX_OUTPUT_CTRL_LANE2 = 32'h00000000;
parameter [31:0] TX_OUTPUT_CTRL_LANE3 = 32'h00000000;
parameter [31:0] TX_OUTPUT_CTRL_LANE4 = 32'h00000000;
parameter [31:0] TX_OUTPUT_CTRL_LANE5 = 32'h00000000;
parameter [31:0] TX_OUTPUT_CTRL_LANE6 = 32'h00000000;
parameter [31:0] TX_OUTPUT_CTRL_LANE7 = 32'h00000000;
parameter [31:0] TX_OUTPUT_EQ_CTRL_LANE0 = 32'h00000000;
parameter [31:0] TX_OUTPUT_EQ_CTRL_LANE1 = 32'h00000000;
parameter [31:0] TX_OUTPUT_EQ_CTRL_LANE2 = 32'h00000000;
parameter [31:0] TX_OUTPUT_EQ_CTRL_LANE3 = 32'h00000000;
parameter [31:0] TX_OUTPUT_EQ_CTRL_LANE4 = 32'h00000000;
parameter [31:0] TX_OUTPUT_EQ_CTRL_LANE5 = 32'h00000000;
parameter [31:0] TX_OUTPUT_EQ_CTRL_LANE6 = 32'h00000000;
parameter [31:0] TX_OUTPUT_EQ_CTRL_LANE7 = 32'h00000000;
parameter [31:0] TX_OUT_LPBK_CTRL_LANE0 = 32'h00000000;
parameter [31:0] TX_OUT_LPBK_CTRL_LANE1 = 32'h00000000;
parameter [31:0] TX_OUT_LPBK_CTRL_LANE2 = 32'h00000000;
parameter [31:0] TX_OUT_LPBK_CTRL_LANE3 = 32'h00000000;
parameter [31:0] TX_OUT_LPBK_CTRL_LANE4 = 32'h00000000;
parameter [31:0] TX_OUT_LPBK_CTRL_LANE5 = 32'h00000000;
parameter [31:0] TX_OUT_LPBK_CTRL_LANE6 = 32'h00000000;
parameter [31:0] TX_OUT_LPBK_CTRL_LANE7 = 32'h00000000;
parameter [31:0] TX_OVERRIDE_CTRL_LANE0 = 32'h00000000;
parameter [31:0] TX_OVERRIDE_CTRL_LANE1 = 32'h00000000;
parameter [31:0] TX_OVERRIDE_CTRL_LANE2 = 32'h00000000;
parameter [31:0] TX_OVERRIDE_CTRL_LANE3 = 32'h00000000;
parameter [31:0] TX_OVERRIDE_CTRL_LANE4 = 32'h00000000;
parameter [31:0] TX_OVERRIDE_CTRL_LANE5 = 32'h00000000;
parameter [31:0] TX_OVERRIDE_CTRL_LANE6 = 32'h00000000;
parameter [31:0] TX_OVERRIDE_CTRL_LANE7 = 32'h00000000;
parameter [31:0] TX_PATTERN_CTRL_LANE0 = 32'h00000000;
parameter [31:0] TX_PATTERN_CTRL_LANE1 = 32'h00000000;
parameter [31:0] TX_PATTERN_CTRL_LANE2 = 32'h00000000;
parameter [31:0] TX_PATTERN_CTRL_LANE3 = 32'h00000000;
parameter [31:0] TX_PATTERN_CTRL_LANE4 = 32'h00000000;
parameter [31:0] TX_PATTERN_CTRL_LANE5 = 32'h00000000;
parameter [31:0] TX_PATTERN_CTRL_LANE6 = 32'h00000000;
parameter [31:0] TX_PATTERN_CTRL_LANE7 = 32'h00000000;
parameter [31:0] TX_PHASE_CTRL_LANE0 = 32'h00000000;
parameter [31:0] TX_PHASE_CTRL_LANE1 = 32'h00000000;
parameter [31:0] TX_PHASE_CTRL_LANE2 = 32'h00000000;
parameter [31:0] TX_PHASE_CTRL_LANE3 = 32'h00000000;
parameter [31:0] TX_PHASE_CTRL_LANE4 = 32'h00000000;
parameter [31:0] TX_PHASE_CTRL_LANE5 = 32'h00000000;
parameter [31:0] TX_PHASE_CTRL_LANE6 = 32'h00000000;
parameter [31:0] TX_PHASE_CTRL_LANE7 = 32'h00000000;
parameter [31:0] TX_REFCLK_SYNC_CTRL_LANE0 = 32'h00000000;
parameter [31:0] TX_REFCLK_SYNC_CTRL_LANE1 = 32'h00000000;
parameter [31:0] TX_REFCLK_SYNC_CTRL_LANE2 = 32'h00000000;
parameter [31:0] TX_REFCLK_SYNC_CTRL_LANE3 = 32'h00000000;
parameter [31:0] TX_REFCLK_SYNC_CTRL_LANE4 = 32'h00000000;
parameter [31:0] TX_REFCLK_SYNC_CTRL_LANE5 = 32'h00000000;
parameter [31:0] TX_REFCLK_SYNC_CTRL_LANE6 = 32'h00000000;
parameter [31:0] TX_REFCLK_SYNC_CTRL_LANE7 = 32'h00000000;
parameter [2:0] TX_SAMPLE_PERIOD_LANE0 = 3'b110;
parameter [2:0] TX_SAMPLE_PERIOD_LANE1 = 3'b110;
parameter [2:0] TX_SAMPLE_PERIOD_LANE2 = 3'b110;
parameter [2:0] TX_SAMPLE_PERIOD_LANE3 = 3'b110;
parameter [2:0] TX_SAMPLE_PERIOD_LANE4 = 3'b110;
parameter [2:0] TX_SAMPLE_PERIOD_LANE5 = 3'b110;
parameter [2:0] TX_SAMPLE_PERIOD_LANE6 = 3'b110;
parameter [2:0] TX_SAMPLE_PERIOD_LANE7 = 3'b110;
parameter [31:0] TX_USER_REG_CTRL_LANE0 = 32'h00000000;
parameter [31:0] TX_USER_REG_CTRL_LANE1 = 32'h00000000;
parameter [31:0] TX_USER_REG_CTRL_LANE2 = 32'h00000000;
parameter [31:0] TX_USER_REG_CTRL_LANE3 = 32'h00000000;
parameter [31:0] TX_USER_REG_CTRL_LANE4 = 32'h00000000;
parameter [31:0] TX_USER_REG_CTRL_LANE5 = 32'h00000000;
parameter [31:0] TX_USER_REG_CTRL_LANE6 = 32'h00000000;
parameter [31:0] TX_USER_REG_CTRL_LANE7 = 32'h00000000;
parameter [31:0] WATCH_DOG_TIMER = 32'h000003E8;
endmodule
//#### END MODULE DEFINITION FOR: GTZE2_OCTAL ####

//#### BEGIN MODULE DEFINITION FOR :IBUF ###
module IBUF (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
parameter CAPACITANCE = "DONT_CARE";
parameter IBUF_DELAY_VALUE = "0";
parameter IBUF_LOW_PWR = "TRUE";
parameter IFD_DELAY_VALUE = "AUTO";
parameter IOSTANDARD = "DEFAULT";
endmodule
//#### END MODULE DEFINITION FOR: IBUF ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS ###
module IBUFDS (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
parameter CAPACITANCE = "DONT_CARE";
parameter DIFF_TERM = "FALSE";
parameter DQS_BIAS = "FALSE";
parameter IBUF_DELAY_VALUE = "0";
parameter IBUF_LOW_PWR = "TRUE";
parameter IFD_DELAY_VALUE = "AUTO";
parameter IOSTANDARD = "DEFAULT";
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_BLVDS_25 ###
module IBUFDS_BLVDS_25 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_BLVDS_25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_DIFF_OUT ###
module IBUFDS_DIFF_OUT (O, OB, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
output OB ;
parameter DIFF_TERM = "FALSE";
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_DIFF_OUT ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_DIFF_OUT_IBUFDISABLE ###
module IBUFDS_DIFF_OUT_IBUFDISABLE (O, OB, I, IB, IBUFDISABLE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
input IBUFDISABLE ;
output O ;
output OB ;
parameter DIFF_TERM = "FALSE";
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
parameter USE_IBUFDISABLE = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_DIFF_OUT_IBUFDISABLE ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_DIFF_OUT_INTERMDISABLE ###
module IBUFDS_DIFF_OUT_INTERMDISABLE (O, OB, I, IB, IBUFDISABLE, INTERMDISABLE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
input IBUFDISABLE ;
input INTERMDISABLE ;
output O ;
output OB ;
parameter DIFF_TERM = "FALSE";
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
parameter USE_IBUFDISABLE = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_DIFF_OUT_INTERMDISABLE ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_DLY_ADJ ###
module IBUFDS_DLY_ADJ (O, I, IB, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
input [2:0] S ;
output O ;
parameter DELAY_OFFSET = "OFF";
parameter DIFF_TERM    = "FALSE";
parameter IOSTANDARD   = "DEFAULT";
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_DLY_ADJ ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_GTE2 ###
module IBUFDS_GTE2 (
  O,
  ODIV2,

  CEB,
  I,
  IB
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CEB ;
input I ;
input IB ;
output O ;
output ODIV2 ;
parameter CLKCM_CFG = "TRUE";
parameter CLKRCV_TRST = "TRUE";
parameter [1:0] CLKSWING_CFG = 2'b11;
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_GTE2 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_GTHE1 ###
module IBUFDS_GTHE1 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_GTHE1 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_GTXE1 ###
module IBUFDS_GTXE1 (O, ODIV2, CEB, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CEB ;
input I ;
input IB ;
output O ;
output ODIV2 ;
parameter CLKCM_CFG = "TRUE";
parameter CLKRCV_TRST = "TRUE";
parameter [9:0] REFCLKOUT_DLY = 10'b0000000000;
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_GTXE1 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_IBUFDISABLE ###
module IBUFDS_IBUFDISABLE (O, I, IB, IBUFDISABLE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
input IBUFDISABLE ;
output O ;
parameter DIFF_TERM = "FALSE";
parameter DQS_BIAS = "FALSE";
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
parameter USE_IBUFDISABLE = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_IBUFDISABLE ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_INTERMDISABLE ###
module IBUFDS_INTERMDISABLE (O, I, IB, IBUFDISABLE, INTERMDISABLE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
input IBUFDISABLE ;
input INTERMDISABLE ;
output O ;
parameter DIFF_TERM = "FALSE";
parameter DQS_BIAS = "FALSE";
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
parameter USE_IBUFDISABLE = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_INTERMDISABLE ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_LDT_25 ###
module IBUFDS_LDT_25 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_LDT_25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_LVDSEXT_25 ###
module IBUFDS_LVDSEXT_25 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_LVDSEXT_25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_LVDSEXT_25_DCI ###
module IBUFDS_LVDSEXT_25_DCI (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_LVDSEXT_25_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_LVDSEXT_33 ###
module IBUFDS_LVDSEXT_33 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_LVDSEXT_33 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_LVDSEXT_33_DCI ###
module IBUFDS_LVDSEXT_33_DCI (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_LVDSEXT_33_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_LVDS_25 ###
module IBUFDS_LVDS_25 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_LVDS_25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_LVDS_25_DCI ###
module IBUFDS_LVDS_25_DCI (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_LVDS_25_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_LVDS_33 ###
module IBUFDS_LVDS_33 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_LVDS_33 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_LVDS_33_DCI ###
module IBUFDS_LVDS_33_DCI (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_LVDS_33_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_LVPECL_25 ###
module IBUFDS_LVPECL_25 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_LVPECL_25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_LVPECL_33 ###
module IBUFDS_LVPECL_33 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_LVPECL_33 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFDS_ULVDS_25 ###
module IBUFDS_ULVDS_25 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFDS_ULVDS_25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG ###
module IBUFG (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
parameter CAPACITANCE = "DONT_CARE";
parameter IBUF_DELAY_VALUE = "0";
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
endmodule
//#### END MODULE DEFINITION FOR: IBUFG ####

//#### BEGIN MODULE DEFINITION FOR :IBUFGDS ###
module IBUFGDS (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
parameter CAPACITANCE = "DONT_CARE";
parameter DIFF_TERM = "FALSE";
parameter IBUF_DELAY_VALUE = "0";
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
endmodule
//#### END MODULE DEFINITION FOR: IBUFGDS ####

//#### BEGIN MODULE DEFINITION FOR :IBUFGDS_BLVDS_25 ###
module IBUFGDS_BLVDS_25 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFGDS_BLVDS_25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFGDS_DIFF_OUT ###
module IBUFGDS_DIFF_OUT (O, OB, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
output OB ;
parameter DIFF_TERM = "FALSE";
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
endmodule
//#### END MODULE DEFINITION FOR: IBUFGDS_DIFF_OUT ####

//#### BEGIN MODULE DEFINITION FOR :IBUFGDS_LDT_25 ###
module IBUFGDS_LDT_25 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFGDS_LDT_25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFGDS_LVDSEXT_25 ###
module IBUFGDS_LVDSEXT_25 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFGDS_LVDSEXT_25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFGDS_LVDSEXT_25_DCI ###
module IBUFGDS_LVDSEXT_25_DCI (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFGDS_LVDSEXT_25_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFGDS_LVDSEXT_33 ###
module IBUFGDS_LVDSEXT_33 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFGDS_LVDSEXT_33 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFGDS_LVDSEXT_33_DCI ###
module IBUFGDS_LVDSEXT_33_DCI (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFGDS_LVDSEXT_33_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFGDS_LVDS_25 ###
module IBUFGDS_LVDS_25 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFGDS_LVDS_25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFGDS_LVDS_25_DCI ###
module IBUFGDS_LVDS_25_DCI (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFGDS_LVDS_25_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFGDS_LVDS_33 ###
module IBUFGDS_LVDS_33 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFGDS_LVDS_33 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFGDS_LVDS_33_DCI ###
module IBUFGDS_LVDS_33_DCI (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFGDS_LVDS_33_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFGDS_LVPECL_25 ###
module IBUFGDS_LVPECL_25 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFGDS_LVPECL_25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFGDS_LVPECL_33 ###
module IBUFGDS_LVPECL_33 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFGDS_LVPECL_33 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFGDS_ULVDS_25 ###
module IBUFGDS_ULVDS_25 (O, I, IB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IB ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFGDS_ULVDS_25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_AGP ###
module IBUFG_AGP (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_AGP ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_CTT ###
module IBUFG_CTT (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_CTT ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_GTL ###
module IBUFG_GTL (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_GTL ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_GTLP ###
module IBUFG_GTLP (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_GTLP ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_GTLP_DCI ###
module IBUFG_GTLP_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_GTLP_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_GTL_DCI ###
module IBUFG_GTL_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_GTL_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_HSTL_I ###
module IBUFG_HSTL_I (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_HSTL_I ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_HSTL_II ###
module IBUFG_HSTL_II (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_HSTL_II ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_HSTL_III ###
module IBUFG_HSTL_III (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_HSTL_III ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_HSTL_III_18 ###
module IBUFG_HSTL_III_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_HSTL_III_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_HSTL_III_DCI ###
module IBUFG_HSTL_III_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_HSTL_III_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_HSTL_III_DCI_18 ###
module IBUFG_HSTL_III_DCI_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_HSTL_III_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_HSTL_II_18 ###
module IBUFG_HSTL_II_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_HSTL_II_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_HSTL_II_DCI ###
module IBUFG_HSTL_II_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_HSTL_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_HSTL_II_DCI_18 ###
module IBUFG_HSTL_II_DCI_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_HSTL_II_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_HSTL_IV ###
module IBUFG_HSTL_IV (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_HSTL_IV ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_HSTL_IV_18 ###
module IBUFG_HSTL_IV_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_HSTL_IV_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_HSTL_IV_DCI ###
module IBUFG_HSTL_IV_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_HSTL_IV_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_HSTL_IV_DCI_18 ###
module IBUFG_HSTL_IV_DCI_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_HSTL_IV_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_HSTL_I_18 ###
module IBUFG_HSTL_I_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_HSTL_I_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_HSTL_I_DCI ###
module IBUFG_HSTL_I_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_HSTL_I_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_HSTL_I_DCI_18 ###
module IBUFG_HSTL_I_DCI_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_HSTL_I_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVCMOS12 ###
module IBUFG_LVCMOS12 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVCMOS12 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVCMOS15 ###
module IBUFG_LVCMOS15 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVCMOS15 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVCMOS18 ###
module IBUFG_LVCMOS18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVCMOS18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVCMOS2 ###
module IBUFG_LVCMOS2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVCMOS2 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVCMOS25 ###
module IBUFG_LVCMOS25 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVCMOS25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVCMOS33 ###
module IBUFG_LVCMOS33 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVCMOS33 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVDCI_15 ###
module IBUFG_LVDCI_15 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVDCI_15 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVDCI_18 ###
module IBUFG_LVDCI_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVDCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVDCI_25 ###
module IBUFG_LVDCI_25 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVDCI_25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVDCI_33 ###
module IBUFG_LVDCI_33 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVDCI_33 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVDCI_DV2_15 ###
module IBUFG_LVDCI_DV2_15 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVDCI_DV2_15 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVDCI_DV2_18 ###
module IBUFG_LVDCI_DV2_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVDCI_DV2_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVDCI_DV2_25 ###
module IBUFG_LVDCI_DV2_25 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVDCI_DV2_25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVDCI_DV2_33 ###
module IBUFG_LVDCI_DV2_33 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVDCI_DV2_33 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVDS ###
module IBUFG_LVDS (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVDS ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVPECL ###
module IBUFG_LVPECL (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVPECL ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_LVTTL ###
module IBUFG_LVTTL (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_LVTTL ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_PCI33_3 ###
module IBUFG_PCI33_3 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_PCI33_3 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_PCI33_5 ###
module IBUFG_PCI33_5 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_PCI33_5 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_PCI66_3 ###
module IBUFG_PCI66_3 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_PCI66_3 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_PCIX ###
module IBUFG_PCIX (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_PCIX ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_PCIX66_3 ###
module IBUFG_PCIX66_3 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_PCIX66_3 ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_SSTL18_I ###
module IBUFG_SSTL18_I (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_SSTL18_I ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_SSTL18_II ###
module IBUFG_SSTL18_II (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_SSTL18_II ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_SSTL18_II_DCI ###
module IBUFG_SSTL18_II_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_SSTL18_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_SSTL18_I_DCI ###
module IBUFG_SSTL18_I_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_SSTL18_I_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_SSTL2_I ###
module IBUFG_SSTL2_I (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_SSTL2_I ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_SSTL2_II ###
module IBUFG_SSTL2_II (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_SSTL2_II ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_SSTL2_II_DCI ###
module IBUFG_SSTL2_II_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_SSTL2_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_SSTL2_I_DCI ###
module IBUFG_SSTL2_I_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_SSTL2_I_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_SSTL3_I ###
module IBUFG_SSTL3_I (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_SSTL3_I ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_SSTL3_II ###
module IBUFG_SSTL3_II (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_SSTL3_II ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_SSTL3_II_DCI ###
module IBUFG_SSTL3_II_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_SSTL3_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUFG_SSTL3_I_DCI ###
module IBUFG_SSTL3_I_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUFG_SSTL3_I_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_AGP ###
module IBUF_AGP (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_AGP ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_CTT ###
module IBUF_CTT (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_CTT ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_DLY_ADJ ###
module IBUF_DLY_ADJ (O, I, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input [2:0] S ;
output O ;
parameter DELAY_OFFSET = "OFF";
parameter IOSTANDARD = "DEFAULT";
endmodule
//#### END MODULE DEFINITION FOR: IBUF_DLY_ADJ ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_GTL ###
module IBUF_GTL (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_GTL ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_GTLP ###
module IBUF_GTLP (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_GTLP ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_GTLP_DCI ###
module IBUF_GTLP_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_GTLP_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_GTL_DCI ###
module IBUF_GTL_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_GTL_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_HSTL_I ###
module IBUF_HSTL_I (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_HSTL_I ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_HSTL_II ###
module IBUF_HSTL_II (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_HSTL_II ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_HSTL_III ###
module IBUF_HSTL_III (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_HSTL_III ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_HSTL_III_18 ###
module IBUF_HSTL_III_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_HSTL_III_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_HSTL_III_DCI ###
module IBUF_HSTL_III_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_HSTL_III_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_HSTL_III_DCI_18 ###
module IBUF_HSTL_III_DCI_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_HSTL_III_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_HSTL_II_18 ###
module IBUF_HSTL_II_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_HSTL_II_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_HSTL_II_DCI ###
module IBUF_HSTL_II_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_HSTL_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_HSTL_II_DCI_18 ###
module IBUF_HSTL_II_DCI_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_HSTL_II_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_HSTL_IV ###
module IBUF_HSTL_IV (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_HSTL_IV ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_HSTL_IV_18 ###
module IBUF_HSTL_IV_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_HSTL_IV_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_HSTL_IV_DCI ###
module IBUF_HSTL_IV_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_HSTL_IV_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_HSTL_IV_DCI_18 ###
module IBUF_HSTL_IV_DCI_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_HSTL_IV_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_HSTL_I_18 ###
module IBUF_HSTL_I_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_HSTL_I_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_HSTL_I_DCI ###
module IBUF_HSTL_I_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_HSTL_I_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_HSTL_I_DCI_18 ###
module IBUF_HSTL_I_DCI_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_HSTL_I_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_IBUFDISABLE ###
module IBUF_IBUFDISABLE (O, I, IBUFDISABLE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IBUFDISABLE ;
output O ;
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
parameter USE_IBUFDISABLE = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: IBUF_IBUFDISABLE ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_INTERMDISABLE ###
module IBUF_INTERMDISABLE (O, I, IBUFDISABLE, INTERMDISABLE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IBUFDISABLE ;
input INTERMDISABLE ;
output O ;
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
parameter USE_IBUFDISABLE = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: IBUF_INTERMDISABLE ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVCMOS12 ###
module IBUF_LVCMOS12 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVCMOS12 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVCMOS15 ###
module IBUF_LVCMOS15 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVCMOS15 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVCMOS18 ###
module IBUF_LVCMOS18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVCMOS18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVCMOS2 ###
module IBUF_LVCMOS2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVCMOS2 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVCMOS25 ###
module IBUF_LVCMOS25 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVCMOS25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVCMOS33 ###
module IBUF_LVCMOS33 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVCMOS33 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVDCI_15 ###
module IBUF_LVDCI_15 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVDCI_15 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVDCI_18 ###
module IBUF_LVDCI_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVDCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVDCI_25 ###
module IBUF_LVDCI_25 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVDCI_25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVDCI_33 ###
module IBUF_LVDCI_33 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVDCI_33 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVDCI_DV2_15 ###
module IBUF_LVDCI_DV2_15 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVDCI_DV2_15 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVDCI_DV2_18 ###
module IBUF_LVDCI_DV2_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVDCI_DV2_18 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVDCI_DV2_25 ###
module IBUF_LVDCI_DV2_25 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVDCI_DV2_25 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVDCI_DV2_33 ###
module IBUF_LVDCI_DV2_33 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVDCI_DV2_33 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVDS ###
module IBUF_LVDS (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVDS ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVPECL ###
module IBUF_LVPECL (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVPECL ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_LVTTL ###
module IBUF_LVTTL (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_LVTTL ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_PCI33_3 ###
module IBUF_PCI33_3 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_PCI33_3 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_PCI33_5 ###
module IBUF_PCI33_5 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_PCI33_5 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_PCI66_3 ###
module IBUF_PCI66_3 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_PCI66_3 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_PCIX ###
module IBUF_PCIX (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_PCIX ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_PCIX66_3 ###
module IBUF_PCIX66_3 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_PCIX66_3 ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_SSTL18_I ###
module IBUF_SSTL18_I (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_SSTL18_I ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_SSTL18_II ###
module IBUF_SSTL18_II (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_SSTL18_II ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_SSTL18_II_DCI ###
module IBUF_SSTL18_II_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_SSTL18_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_SSTL18_I_DCI ###
module IBUF_SSTL18_I_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_SSTL18_I_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_SSTL2_I ###
module IBUF_SSTL2_I (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_SSTL2_I ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_SSTL2_II ###
module IBUF_SSTL2_II (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_SSTL2_II ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_SSTL2_II_DCI ###
module IBUF_SSTL2_II_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_SSTL2_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_SSTL2_I_DCI ###
module IBUF_SSTL2_I_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_SSTL2_I_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_SSTL3_I ###
module IBUF_SSTL3_I (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_SSTL3_I ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_SSTL3_II ###
module IBUF_SSTL3_II (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_SSTL3_II ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_SSTL3_II_DCI ###
module IBUF_SSTL3_II_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_SSTL3_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IBUF_SSTL3_I_DCI ###
module IBUF_SSTL3_I_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: IBUF_SSTL3_I_DCI ####

//#### BEGIN MODULE DEFINITION FOR :ICAPE2 ###
module ICAPE2 (
  O,
  CLK,
  CSIB,
  I,
  RDWRB
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLK ;
input CSIB ;
input RDWRB ;
input [31:0] I ;
output [31:0] O ;
parameter [31:0] DEVICE_ID = 32'h03651093;
parameter ICAP_WIDTH = "X32";
parameter SIM_CFG_FILE_NAME = "NONE";
endmodule
//#### END MODULE DEFINITION FOR: ICAPE2 ####

//#### BEGIN MODULE DEFINITION FOR :ICAP_SPARTAN3A ###
module ICAP_SPARTAN3A (BUSY, O, CE, CLK, I, WRITE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CE ;
input CLK ;
input WRITE ;
input [7:0] I ;
output BUSY ;
output [7:0] O ;
endmodule
//#### END MODULE DEFINITION FOR: ICAP_SPARTAN3A ####

//#### BEGIN MODULE DEFINITION FOR :ICAP_SPARTAN6 ###
module ICAP_SPARTAN6 (
  BUSY,
  O,
  CE,
  CLK,
  I,
  WRITE
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLK ;
input CE ;
input WRITE ;
input [15:0] I ;
output BUSY ;
output [15:0] O ;
parameter DEVICE_ID = 32'h04000093;
parameter SIM_CFG_FILE_NAME = "NONE";
endmodule
//#### END MODULE DEFINITION FOR: ICAP_SPARTAN6 ####

//#### BEGIN MODULE DEFINITION FOR :ICAP_VIRTEX4 ###
module ICAP_VIRTEX4 (BUSY, O, CE, CLK, I, WRITE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CE ;
input CLK ;
input WRITE ;
input [31:0] I ;
output BUSY ;
output [31:0] O ;
parameter ICAP_WIDTH = "X8";
endmodule
//#### END MODULE DEFINITION FOR: ICAP_VIRTEX4 ####

//#### BEGIN MODULE DEFINITION FOR :ICAP_VIRTEX5 ###
module ICAP_VIRTEX5 (
	BUSY,
	O,
	CE,
	CLK,
	I,
	WRITE
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CE ;
input CLK ;
input WRITE ;
input [31:0] I ;
output BUSY ;
output [31:0] O ;
parameter ICAP_WIDTH = "X8";
endmodule
//#### END MODULE DEFINITION FOR: ICAP_VIRTEX5 ####

//#### BEGIN MODULE DEFINITION FOR :ICAP_VIRTEX6 ###
module ICAP_VIRTEX6 (
  BUSY,
  O,
  CLK,
  CSB,
  I,
  RDWRB
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLK ;
input CSB ;
input RDWRB ;
input [31:0] I ;
output BUSY ;
output [31:0] O ;
parameter [31:0] DEVICE_ID = 32'h04244093;
parameter ICAP_WIDTH = "X8";
parameter SIM_CFG_FILE_NAME = "NONE";
endmodule
//#### END MODULE DEFINITION FOR: ICAP_VIRTEX6 ####

//#### BEGIN MODULE DEFINITION FOR :IDDR ###
module IDDR (Q1, Q2, C, CE, D, R, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input D ;
input R ;
input S ;
output Q1 ;
output Q2 ;
parameter DDR_CLK_EDGE = "OPPOSITE_EDGE";
parameter INIT_Q1 = 1'b0;
parameter INIT_Q2 = 1'b0;
parameter SRTYPE = "SYNC";
endmodule
//#### END MODULE DEFINITION FOR: IDDR ####

//#### BEGIN MODULE DEFINITION FOR :IDDR2 ###
module IDDR2 (Q0, Q1, C0, C1, CE, D, R, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C0 ;
input C1 ;
input CE ;
input D ;
input R ;
input S ;
output Q0 ;
output Q1 ;
parameter DDR_ALIGNMENT = "NONE";
parameter INIT_Q0 = 1'b0;
parameter INIT_Q1 = 1'b0;
parameter SRTYPE = "SYNC";
endmodule
//#### END MODULE DEFINITION FOR: IDDR2 ####

//#### BEGIN MODULE DEFINITION FOR :IDDR_2CLK ###
module IDDR_2CLK (Q1, Q2, C, CB, CE, D, R, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CB ;
input CE ;
input D ;
input R ;
input S ;
output Q1 ;
output Q2 ;
parameter DDR_CLK_EDGE = "OPPOSITE_EDGE";
parameter INIT_Q1 = 1'b0;
parameter INIT_Q2 = 1'b0;
parameter SRTYPE = "SYNC";
endmodule
//#### END MODULE DEFINITION FOR: IDDR_2CLK ####

//#### BEGIN MODULE DEFINITION FOR :IDELAY ###
module IDELAY (O, C, CE, I, INC, RST) /* synthesis syn_black_box  syn_lib_cell=1
 .noprune=1
 */;
input C ;
input CE ;
input I ;
input INC ;
input RST ;
output O ;
parameter IOBDELAY_TYPE = "DEFAULT";
parameter IOBDELAY_VALUE = 0;
endmodule
//#### END MODULE DEFINITION FOR: IDELAY ####

//#### BEGIN MODULE DEFINITION FOR :IDELAYCTRL ###
module IDELAYCTRL (RDY, REFCLK, RST) /* synthesis syn_black_box  syn_lib_cell=1
 .noprune=1
 */;
input REFCLK ;
input RST ;
output RDY ;
endmodule
//#### END MODULE DEFINITION FOR: IDELAYCTRL ####

//#### BEGIN MODULE DEFINITION FOR :IDELAYE2 ###
module IDELAYE2 (CNTVALUEOUT, DATAOUT, C, CE, CINVCTRL, CNTVALUEIN, DATAIN, IDATAIN, INC, LD, LDPIPEEN, REGRST) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input CINVCTRL ;
input [4:0] CNTVALUEIN ;
input DATAIN ;
input IDATAIN ;
input INC ;
input LD ;
input LDPIPEEN ;
input REGRST ;
output [4:0] CNTVALUEOUT ;
output DATAOUT ;
parameter CINVCTRL_SEL = "FALSE";
parameter DELAY_SRC = "IDATAIN";
parameter HIGH_PERFORMANCE_MODE    = "FALSE";
parameter IDELAY_TYPE  = "FIXED";
parameter IDELAY_VALUE = 0;
parameter PIPE_SEL = "FALSE";
parameter REFCLK_FREQUENCY = 200.0;
parameter SIGNAL_PATTERN    = "DATA";
endmodule
//#### END MODULE DEFINITION FOR: IDELAYE2 ####

//#### BEGIN MODULE DEFINITION FOR :IDELAYE2_FINEDELAY ###
module IDELAYE2_FINEDELAY (
  CNTVALUEOUT,
  DATAOUT,

  C,
  CE,
  CINVCTRL,
  CNTVALUEIN,
  DATAIN,
  IDATAIN,
  IFDLY,
  INC,
  LD,
  LDPIPEEN,
  REGRST
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input CINVCTRL ;
input [4:0] CNTVALUEIN ;
input DATAIN ;
input IDATAIN ;
input [2:0] IFDLY ;
input INC ;
input LD ;
input LDPIPEEN ;
input REGRST ;
output [4:0] CNTVALUEOUT ;
output DATAOUT ;
parameter CINVCTRL_SEL = "FALSE";
parameter DELAY_SRC = "IDATAIN";
parameter FINEDELAY = "BYPASS";
parameter HIGH_PERFORMANCE_MODE    = "FALSE";
parameter IDELAY_TYPE  = "FIXED";
parameter IDELAY_VALUE = 0;
parameter PIPE_SEL = "FALSE";
parameter REFCLK_FREQUENCY = 200.0;
parameter SIGNAL_PATTERN    = "DATA";
endmodule
//#### END MODULE DEFINITION FOR: IDELAYE2_FINEDELAY ####

//#### BEGIN MODULE DEFINITION FOR :IFDDRCPE ###
module IFDDRCPE (Q0, Q1, C0, C1, CE, CLR, D, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C0 ;
input C1 ;
input CE ;
input CLR ;
input D ;
input PRE ;
output Q0 ;
output Q1 ;
endmodule
//#### END MODULE DEFINITION FOR: IFDDRCPE ####

//#### BEGIN MODULE DEFINITION FOR :IFDDRRSE ###
module IFDDRRSE (Q0, Q1, C0, C1, CE, D, R, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C0 ;
input C1 ;
input CE ;
input D ;
input R ;
input S ;
output Q0 ;
output Q1 ;
endmodule
//#### END MODULE DEFINITION FOR: IFDDRRSE ####

//#### BEGIN MODULE DEFINITION FOR :INV ###
module INV (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: INV ####

//#### BEGIN MODULE DEFINITION FOR :IN_FIFO ###
module IN_FIFO (
  ALMOSTEMPTY,
  ALMOSTFULL,
  EMPTY,
  FULL,
  Q0,
  Q1,
  Q2,
  Q3,
  Q4,
  Q5,
  Q6,
  Q7,
  Q8,
  Q9,

  D0,
  D1,
  D2,
  D3,
  D4,
  D5,
  D6,
  D7,
  D8,
  D9,
  RDCLK,
  RDEN,
  RESET,
  WRCLK,
  WREN
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input RDCLK ;
input RDEN ;
input RESET ;
input WRCLK ;
input WREN ;
input [3:0] D0 ;
input [3:0] D1 ;
input [3:0] D2 ;
input [3:0] D3 ;
input [3:0] D4 ;
input [3:0] D7 ;
input [3:0] D8 ;
input [3:0] D9 ;
input [7:0] D5 ;
input [7:0] D6 ;
output ALMOSTEMPTY ;
output ALMOSTFULL ;
output EMPTY ;
output FULL ;
output [7:0] Q0 ;
output [7:0] Q1 ;
output [7:0] Q2 ;
output [7:0] Q3 ;
output [7:0] Q4 ;
output [7:0] Q5 ;
output [7:0] Q6 ;
output [7:0] Q7 ;
output [7:0] Q8 ;
output [7:0] Q9 ;
parameter ALMOST_EMPTY_VALUE = 1;
parameter ALMOST_FULL_VALUE = 1;
parameter ARRAY_MODE = "ARRAY_MODE_4_X_8";
parameter SYNCHRONOUS_MODE = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: IN_FIFO ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF ###
module IOBUF (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
parameter CAPACITANCE = "DONT_CARE";
parameter DRIVE = 12;
parameter IBUF_DELAY_VALUE = "0";
parameter IBUF_LOW_PWR = "TRUE";
parameter IFD_DELAY_VALUE = "AUTO";
parameter IOSTANDARD = "DEFAULT";
parameter SLEW = "SLOW";
endmodule
//#### END MODULE DEFINITION FOR: IOBUF ####

//#### BEGIN MODULE DEFINITION FOR :IOBUFDS ###
module IOBUFDS (O, IO, IOB, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
inout IOB ;
parameter CAPACITANCE = "DONT_CARE";
parameter DIFF_TERM = "FALSE";
parameter DQS_BIAS = "FALSE";
parameter IBUF_DELAY_VALUE = "0";
parameter IBUF_LOW_PWR = "TRUE";
parameter IFD_DELAY_VALUE = "AUTO";
parameter IOSTANDARD = "DEFAULT";
parameter SLEW = "SLOW";
endmodule
//#### END MODULE DEFINITION FOR: IOBUFDS ####

//#### BEGIN MODULE DEFINITION FOR :IOBUFDS_BLVDS_25 ###
module IOBUFDS_BLVDS_25 (O, IO, IOB, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
inout IOB ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUFDS_BLVDS_25 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUFDS_DCIEN ###
module IOBUFDS_DCIEN (O, IO, IOB, DCITERMDISABLE, I, IBUFDISABLE, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input DCITERMDISABLE ;
input I ;
input IBUFDISABLE ;
input T ;
output O ;
inout IO ;
inout IOB ;
parameter DIFF_TERM = "FALSE";
parameter DQS_BIAS = "FALSE";
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
parameter SLEW = "SLOW";
parameter USE_IBUFDISABLE = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: IOBUFDS_DCIEN ####

//#### BEGIN MODULE DEFINITION FOR :IOBUFDS_DIFF_OUT ###
module IOBUFDS_DIFF_OUT (O, OB, IO, IOB, I, TM, TS) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input TM ;
input TS ;
output O ;
output OB ;
inout IO ;
inout IOB ;
parameter DIFF_TERM = "FALSE";
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
endmodule
//#### END MODULE DEFINITION FOR: IOBUFDS_DIFF_OUT ####

//#### BEGIN MODULE DEFINITION FOR :IOBUFDS_DIFF_OUT_DCIEN ###
module IOBUFDS_DIFF_OUT_DCIEN (O, OB, IO, IOB, DCITERMDISABLE, I, IBUFDISABLE, TM, TS) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input DCITERMDISABLE ;
input I ;
input IBUFDISABLE ;
input TM ;
input TS ;
output O ;
output OB ;
inout IO ;
inout IOB ;
parameter DIFF_TERM = "FALSE";
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
parameter USE_IBUFDISABLE = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: IOBUFDS_DIFF_OUT_DCIEN ####

//#### BEGIN MODULE DEFINITION FOR :IOBUFDS_DIFF_OUT_INTERMDISABLE ###
module IOBUFDS_DIFF_OUT_INTERMDISABLE (O, OB, IO, IOB, I, IBUFDISABLE, INTERMDISABLE, TM, TS) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IBUFDISABLE ;
input INTERMDISABLE ;
input TM ;
input TS ;
output O ;
output OB ;
inout IO ;
inout IOB ;
parameter DIFF_TERM = "FALSE";
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
parameter USE_IBUFDISABLE = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: IOBUFDS_DIFF_OUT_INTERMDISABLE ####

//#### BEGIN MODULE DEFINITION FOR :IOBUFDS_INTERMDISABLE ###
module IOBUFDS_INTERMDISABLE (O, IO, IOB, I, IBUFDISABLE, INTERMDISABLE, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IBUFDISABLE ;
input INTERMDISABLE ;
input T ;
output O ;
inout IO ;
inout IOB ;
parameter DIFF_TERM = "FALSE";
parameter DQS_BIAS = "FALSE";
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
parameter SLEW = "SLOW";
parameter USE_IBUFDISABLE = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: IOBUFDS_INTERMDISABLE ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_AGP ###
module IOBUF_AGP (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_AGP ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_CTT ###
module IOBUF_CTT (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_CTT ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_DCIEN ###
module IOBUF_DCIEN (O, IO, DCITERMDISABLE, I, IBUFDISABLE, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input DCITERMDISABLE ;
input I ;
input IBUFDISABLE ;
input T ;
output O ;
inout IO ;
parameter DRIVE = 12;
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
parameter SLEW = "SLOW";
parameter USE_IBUFDISABLE = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_DCIEN ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_F_12 ###
module IOBUF_F_12 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_F_16 ###
module IOBUF_F_16 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_F_2 ###
module IOBUF_F_2 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_F_24 ###
module IOBUF_F_24 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_F_24 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_F_4 ###
module IOBUF_F_4 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_F_6 ###
module IOBUF_F_6 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_F_8 ###
module IOBUF_F_8 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_GTL ###
module IOBUF_GTL (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_GTL ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_GTLP ###
module IOBUF_GTLP (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_GTLP ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_GTLP_DCI ###
module IOBUF_GTLP_DCI (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_GTLP_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_GTL_DCI ###
module IOBUF_GTL_DCI (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_GTL_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_HSTL_I ###
module IOBUF_HSTL_I (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_HSTL_I ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_HSTL_II ###
module IOBUF_HSTL_II (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_HSTL_II ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_HSTL_III ###
module IOBUF_HSTL_III (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_HSTL_III ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_HSTL_III_18 ###
module IOBUF_HSTL_III_18 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_HSTL_III_18 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_HSTL_II_18 ###
module IOBUF_HSTL_II_18 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_HSTL_II_18 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_HSTL_II_DCI ###
module IOBUF_HSTL_II_DCI (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_HSTL_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_HSTL_II_DCI_18 ###
module IOBUF_HSTL_II_DCI_18 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_HSTL_II_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_HSTL_IV ###
module IOBUF_HSTL_IV (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_HSTL_IV ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_HSTL_IV_18 ###
module IOBUF_HSTL_IV_18 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_HSTL_IV_18 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_HSTL_IV_DCI ###
module IOBUF_HSTL_IV_DCI (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_HSTL_IV_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_HSTL_IV_DCI_18 ###
module IOBUF_HSTL_IV_DCI_18 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_HSTL_IV_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_HSTL_I_18 ###
module IOBUF_HSTL_I_18 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_HSTL_I_18 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_INTERMDISABLE ###
module IOBUF_INTERMDISABLE (O, IO, I, IBUFDISABLE, INTERMDISABLE, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input IBUFDISABLE ;
input INTERMDISABLE ;
input T ;
output O ;
inout IO ;
parameter DRIVE = 12;
parameter IBUF_LOW_PWR = "TRUE";
parameter IOSTANDARD = "DEFAULT";
parameter SLEW = "SLOW";
parameter USE_IBUFDISABLE = "TRUE";
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_INTERMDISABLE ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS12 ###
module IOBUF_LVCMOS12 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS12 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS12_F_2 ###
module IOBUF_LVCMOS12_F_2 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS12_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS12_F_4 ###
module IOBUF_LVCMOS12_F_4 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS12_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS12_F_6 ###
module IOBUF_LVCMOS12_F_6 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS12_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS12_F_8 ###
module IOBUF_LVCMOS12_F_8 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS12_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS12_S_2 ###
module IOBUF_LVCMOS12_S_2 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS12_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS12_S_4 ###
module IOBUF_LVCMOS12_S_4 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS12_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS12_S_6 ###
module IOBUF_LVCMOS12_S_6 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS12_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS12_S_8 ###
module IOBUF_LVCMOS12_S_8 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS12_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS15 ###
module IOBUF_LVCMOS15 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS15 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS15_F_12 ###
module IOBUF_LVCMOS15_F_12 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS15_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS15_F_16 ###
module IOBUF_LVCMOS15_F_16 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS15_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS15_F_2 ###
module IOBUF_LVCMOS15_F_2 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS15_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS15_F_4 ###
module IOBUF_LVCMOS15_F_4 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS15_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS15_F_6 ###
module IOBUF_LVCMOS15_F_6 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS15_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS15_F_8 ###
module IOBUF_LVCMOS15_F_8 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS15_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS15_S_12 ###
module IOBUF_LVCMOS15_S_12 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS15_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS15_S_16 ###
module IOBUF_LVCMOS15_S_16 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS15_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS15_S_2 ###
module IOBUF_LVCMOS15_S_2 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS15_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS15_S_4 ###
module IOBUF_LVCMOS15_S_4 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS15_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS15_S_6 ###
module IOBUF_LVCMOS15_S_6 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS15_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS15_S_8 ###
module IOBUF_LVCMOS15_S_8 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS15_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS18 ###
module IOBUF_LVCMOS18 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS18 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS18_F_12 ###
module IOBUF_LVCMOS18_F_12 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS18_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS18_F_16 ###
module IOBUF_LVCMOS18_F_16 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS18_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS18_F_2 ###
module IOBUF_LVCMOS18_F_2 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS18_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS18_F_4 ###
module IOBUF_LVCMOS18_F_4 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS18_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS18_F_6 ###
module IOBUF_LVCMOS18_F_6 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS18_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS18_F_8 ###
module IOBUF_LVCMOS18_F_8 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS18_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS18_S_12 ###
module IOBUF_LVCMOS18_S_12 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS18_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS18_S_16 ###
module IOBUF_LVCMOS18_S_16 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS18_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS18_S_2 ###
module IOBUF_LVCMOS18_S_2 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS18_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS18_S_4 ###
module IOBUF_LVCMOS18_S_4 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS18_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS18_S_6 ###
module IOBUF_LVCMOS18_S_6 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS18_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS18_S_8 ###
module IOBUF_LVCMOS18_S_8 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS18_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS2 ###
module IOBUF_LVCMOS2 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS2 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS25 ###
module IOBUF_LVCMOS25 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS25 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS25_F_12 ###
module IOBUF_LVCMOS25_F_12 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS25_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS25_F_16 ###
module IOBUF_LVCMOS25_F_16 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS25_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS25_F_2 ###
module IOBUF_LVCMOS25_F_2 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS25_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS25_F_24 ###
module IOBUF_LVCMOS25_F_24 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS25_F_24 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS25_F_4 ###
module IOBUF_LVCMOS25_F_4 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS25_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS25_F_6 ###
module IOBUF_LVCMOS25_F_6 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS25_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS25_F_8 ###
module IOBUF_LVCMOS25_F_8 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS25_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS25_S_12 ###
module IOBUF_LVCMOS25_S_12 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS25_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS25_S_16 ###
module IOBUF_LVCMOS25_S_16 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS25_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS25_S_2 ###
module IOBUF_LVCMOS25_S_2 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS25_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS25_S_24 ###
module IOBUF_LVCMOS25_S_24 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS25_S_24 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS25_S_4 ###
module IOBUF_LVCMOS25_S_4 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS25_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS25_S_6 ###
module IOBUF_LVCMOS25_S_6 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS25_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS25_S_8 ###
module IOBUF_LVCMOS25_S_8 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS25_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS33 ###
module IOBUF_LVCMOS33 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS33 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS33_F_12 ###
module IOBUF_LVCMOS33_F_12 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS33_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS33_F_16 ###
module IOBUF_LVCMOS33_F_16 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS33_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS33_F_2 ###
module IOBUF_LVCMOS33_F_2 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS33_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS33_F_24 ###
module IOBUF_LVCMOS33_F_24 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS33_F_24 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS33_F_4 ###
module IOBUF_LVCMOS33_F_4 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS33_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS33_F_6 ###
module IOBUF_LVCMOS33_F_6 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS33_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS33_F_8 ###
module IOBUF_LVCMOS33_F_8 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS33_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS33_S_12 ###
module IOBUF_LVCMOS33_S_12 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS33_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS33_S_16 ###
module IOBUF_LVCMOS33_S_16 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS33_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS33_S_2 ###
module IOBUF_LVCMOS33_S_2 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS33_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS33_S_24 ###
module IOBUF_LVCMOS33_S_24 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS33_S_24 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS33_S_4 ###
module IOBUF_LVCMOS33_S_4 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS33_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS33_S_6 ###
module IOBUF_LVCMOS33_S_6 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS33_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVCMOS33_S_8 ###
module IOBUF_LVCMOS33_S_8 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVCMOS33_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVDCI_15 ###
module IOBUF_LVDCI_15 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVDCI_15 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVDCI_18 ###
module IOBUF_LVDCI_18 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVDCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVDCI_25 ###
module IOBUF_LVDCI_25 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVDCI_25 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVDCI_33 ###
module IOBUF_LVDCI_33 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVDCI_33 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVDCI_DV2_15 ###
module IOBUF_LVDCI_DV2_15 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVDCI_DV2_15 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVDCI_DV2_18 ###
module IOBUF_LVDCI_DV2_18 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVDCI_DV2_18 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVDCI_DV2_25 ###
module IOBUF_LVDCI_DV2_25 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVDCI_DV2_25 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVDCI_DV2_33 ###
module IOBUF_LVDCI_DV2_33 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVDCI_DV2_33 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVDS ###
module IOBUF_LVDS (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVDS ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVPECL ###
module IOBUF_LVPECL (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVPECL ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVTTL ###
module IOBUF_LVTTL (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVTTL ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVTTL_F_12 ###
module IOBUF_LVTTL_F_12 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVTTL_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVTTL_F_16 ###
module IOBUF_LVTTL_F_16 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVTTL_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVTTL_F_2 ###
module IOBUF_LVTTL_F_2 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVTTL_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVTTL_F_24 ###
module IOBUF_LVTTL_F_24 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVTTL_F_24 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVTTL_F_4 ###
module IOBUF_LVTTL_F_4 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVTTL_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVTTL_F_6 ###
module IOBUF_LVTTL_F_6 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVTTL_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVTTL_F_8 ###
module IOBUF_LVTTL_F_8 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVTTL_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVTTL_S_12 ###
module IOBUF_LVTTL_S_12 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVTTL_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVTTL_S_16 ###
module IOBUF_LVTTL_S_16 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVTTL_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVTTL_S_2 ###
module IOBUF_LVTTL_S_2 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVTTL_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVTTL_S_24 ###
module IOBUF_LVTTL_S_24 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVTTL_S_24 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVTTL_S_4 ###
module IOBUF_LVTTL_S_4 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVTTL_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVTTL_S_6 ###
module IOBUF_LVTTL_S_6 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVTTL_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_LVTTL_S_8 ###
module IOBUF_LVTTL_S_8 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_LVTTL_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_PCI33_3 ###
module IOBUF_PCI33_3 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_PCI33_3 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_PCI33_5 ###
module IOBUF_PCI33_5 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_PCI33_5 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_PCI66_3 ###
module IOBUF_PCI66_3 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_PCI66_3 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_PCIX ###
module IOBUF_PCIX (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_PCIX ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_PCIX66_3 ###
module IOBUF_PCIX66_3 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_PCIX66_3 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_SSTL18_I ###
module IOBUF_SSTL18_I (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_SSTL18_I ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_SSTL18_II ###
module IOBUF_SSTL18_II (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_SSTL18_II ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_SSTL18_II_DCI ###
module IOBUF_SSTL18_II_DCI (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_SSTL18_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_SSTL2_I ###
module IOBUF_SSTL2_I (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_SSTL2_I ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_SSTL2_II ###
module IOBUF_SSTL2_II (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_SSTL2_II ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_SSTL2_II_DCI ###
module IOBUF_SSTL2_II_DCI (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_SSTL2_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_SSTL3_I ###
module IOBUF_SSTL3_I (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_SSTL3_I ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_SSTL3_II ###
module IOBUF_SSTL3_II (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_SSTL3_II ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_SSTL3_II_DCI ###
module IOBUF_SSTL3_II_DCI (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_SSTL3_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_S_12 ###
module IOBUF_S_12 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_S_16 ###
module IOBUF_S_16 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_S_2 ###
module IOBUF_S_2 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_S_24 ###
module IOBUF_S_24 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_S_24 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_S_4 ###
module IOBUF_S_4 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_S_6 ###
module IOBUF_S_6 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :IOBUF_S_8 ###
module IOBUF_S_8 (O, IO, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O ;
inout IO ;
endmodule
//#### END MODULE DEFINITION FOR: IOBUF_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :IODELAY ###
module IODELAY (DATAOUT, C, CE, DATAIN, IDATAIN, INC, ODATAIN, RST, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input DATAIN ;
input IDATAIN ;
input INC ;
input ODATAIN ;
input RST ;
input T ;
output DATAOUT ;
parameter DELAY_SRC    = "I";
parameter HIGH_PERFORMANCE_MODE    = "TRUE";
parameter IDELAY_TYPE  = "DEFAULT";
parameter IDELAY_VALUE = 0;
parameter ODELAY_VALUE = 0;
parameter REFCLK_FREQUENCY = 200.0;
parameter SIGNAL_PATTERN    = "DATA";
endmodule
//#### END MODULE DEFINITION FOR: IODELAY ####

//#### BEGIN MODULE DEFINITION FOR :IODELAY2 ###
module IODELAY2 (
  BUSY,
  DATAOUT,
  DATAOUT2,
  DOUT,
  TOUT,
  CAL,
  CE,
  CLK,
  IDATAIN,
  INC,
  IOCLK0,
  IOCLK1,
  ODATAIN,
  RST,
  T
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CAL ;
input CE ;
input CLK ;
input IDATAIN ;
input INC ;
input IOCLK0 ;
input IOCLK1 ;
input ODATAIN ;
input RST ;
input T ;
output BUSY ;
output DATAOUT2 ;
output DATAOUT ;
output DOUT ;
output TOUT ;
parameter COUNTER_WRAPAROUND = "WRAPAROUND";
parameter DATA_RATE = "SDR";
parameter DELAY_SRC = "IO";
parameter IDELAY2_VALUE = 0;
parameter IDELAY_MODE = "NORMAL";
parameter IDELAY_TYPE = "DEFAULT";
parameter IDELAY_VALUE = 0;
parameter ODELAY_VALUE = 0;
parameter SERDES_MODE = "NONE";
parameter SIM_TAPDELAY_VALUE = 75;
endmodule
//#### END MODULE DEFINITION FOR: IODELAY2 ####

//#### BEGIN MODULE DEFINITION FOR :IODELAYE1 ###
module IODELAYE1 (CNTVALUEOUT, DATAOUT, C, CE, CINVCTRL, CLKIN, CNTVALUEIN, DATAIN, IDATAIN, INC, ODATAIN, RST, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input CINVCTRL ;
input CLKIN ;
input [4:0] CNTVALUEIN ;
input DATAIN ;
input IDATAIN ;
input INC ;
input ODATAIN ;
input RST ;
input T ;
output [4:0] CNTVALUEOUT ;
output DATAOUT ;
parameter CINVCTRL_SEL = "FALSE";
parameter DELAY_SRC    = "I";
parameter HIGH_PERFORMANCE_MODE    = "FALSE";
parameter IDELAY_TYPE  = "DEFAULT";
parameter IDELAY_VALUE = 0;
parameter ODELAY_TYPE  = "FIXED";
parameter ODELAY_VALUE = 0;
parameter REFCLK_FREQUENCY = 200.0;
parameter SIGNAL_PATTERN    = "DATA";
endmodule
//#### END MODULE DEFINITION FOR: IODELAYE1 ####

//#### BEGIN MODULE DEFINITION FOR :IODRP2 ###
module IODRP2 (
  DATAOUT,
  DATAOUT2,
  DOUT,
  SDO,
  TOUT,
  ADD,
  BKST,
  CLK,
  CS,
  IDATAIN,
  IOCLK0,
  IOCLK1,
  ODATAIN,
  SDI,
  T
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input ADD ;
input BKST ;
input CLK ;
input CS ;
input IDATAIN ;
input IOCLK0 ;
input IOCLK1 ;
input ODATAIN ;
input SDI ;
input T ;
output DATAOUT2 ;
output DATAOUT ;
output DOUT ;
output SDO ;
output TOUT ;
parameter DATA_RATE = "SDR";
parameter SIM_TAPDELAY_VALUE = 75;
endmodule
//#### END MODULE DEFINITION FOR: IODRP2 ####

//#### BEGIN MODULE DEFINITION FOR :IODRP2_MCB ###
module IODRP2_MCB (
  AUXSDO,
  DATAOUT,
  DATAOUT2,
  DOUT,
  DQSOUTN,
  DQSOUTP,
  SDO,
  TOUT,
  ADD,
  AUXADDR,
  AUXSDOIN,
  BKST,
  CLK,
  CS,
  IDATAIN,
  IOCLK0,
  IOCLK1,
  MEMUPDATE,
  ODATAIN,
  SDI,
  T
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input ADD ;
input AUXSDOIN ;
input BKST ;
input CLK ;
input CS ;
input IDATAIN ;
input IOCLK0 ;
input IOCLK1 ;
input MEMUPDATE ;
input ODATAIN ;
input SDI ;
input T ;
input [4:0] AUXADDR ;
output AUXSDO ;
output DATAOUT2 ;
output DATAOUT ;
output DOUT ;
output DQSOUTN ;
output DQSOUTP ;
output SDO ;
output TOUT ;
parameter DATA_RATE = "SDR";
parameter IDELAY_VALUE = 0;
parameter MCB_ADDRESS = 0;
parameter ODELAY_VALUE = 0;
parameter SERDES_MODE = "NONE";
parameter SIM_TAPDELAY_VALUE = 75;
endmodule
//#### END MODULE DEFINITION FOR: IODRP2_MCB ####

//#### BEGIN MODULE DEFINITION FOR :ISERDES ###
module ISERDES (O, Q1, Q2, Q3, Q4, Q5, Q6, SHIFTOUT1, SHIFTOUT2,
		  BITSLIP, CE1, CE2, CLK, CLKDIV, D, DLYCE, DLYINC, DLYRST, OCLK, REV, SHIFTIN1, SHIFTIN2, SR) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input BITSLIP ;
input CE1 ;
input CE2 ;
input CLK ;
input CLKDIV ;
input D ;
input DLYCE ;
input DLYINC ;
input DLYRST ;
input OCLK ;
input REV ;
input SHIFTIN1 ;
input SHIFTIN2 ;
input SR ;
output O ;
output Q1 ;
output Q2 ;
output Q3 ;
output Q4 ;
output Q5 ;
output Q6 ;
output SHIFTOUT1 ;
output SHIFTOUT2 ;
parameter BITSLIP_ENABLE = "FALSE";
parameter DATA_RATE = "DDR";
parameter DATA_WIDTH = 4;
parameter INIT_Q1 = 1'b0;
parameter INIT_Q2 = 1'b0;
parameter INIT_Q3 = 1'b0;
parameter INIT_Q4 = 1'b0;
parameter INTERFACE_TYPE = "MEMORY";
parameter IOBDELAY = "NONE";
parameter IOBDELAY_TYPE = "DEFAULT";
parameter IOBDELAY_VALUE = 0;
parameter NUM_CE = 2;
parameter SERDES_MODE = "MASTER";
parameter SRVAL_Q1 = 1'b0;
parameter SRVAL_Q2 = 1'b0;
parameter SRVAL_Q3 = 1'b0;
parameter SRVAL_Q4 = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: ISERDES ####

//#### BEGIN MODULE DEFINITION FOR :ISERDES2 ###
module ISERDES2 (
  CFB0,
  CFB1,
  DFB,
  FABRICOUT,
  INCDEC,
  Q1,
  Q2,
  Q3,
  Q4,
  SHIFTOUT,
  VALID,
  BITSLIP,
  CE0,
  CLK0,
  CLK1,
  CLKDIV,
  D,
  IOCE,
  RST,
  SHIFTIN
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input BITSLIP ;
input CE0 ;
input CLK0 ;
input CLK1 ;
input CLKDIV ;
input D ;
input IOCE ;
input RST ;
input SHIFTIN ;
output CFB0 ;
output CFB1 ;
output DFB ;
output FABRICOUT ;
output INCDEC ;
output Q1 ;
output Q2 ;
output Q3 ;
output Q4 ;
output SHIFTOUT ;
output VALID ;
parameter BITSLIP_ENABLE = "FALSE";
parameter DATA_RATE = "SDR";
parameter DATA_WIDTH = 1;
parameter INTERFACE_TYPE = "NETWORKING";
parameter SERDES_MODE = "NONE";
endmodule
//#### END MODULE DEFINITION FOR: ISERDES2 ####

//#### BEGIN MODULE DEFINITION FOR :ISERDESE1 ###
module ISERDESE1 (O, Q1, Q2, Q3, Q4, Q5, Q6, SHIFTOUT1, SHIFTOUT2,
                  BITSLIP, CE1, CE2, CLK, CLKB, CLKDIV, D, DDLY, DYNCLKDIVSEL, DYNCLKSEL, OCLK, OFB, RST, SHIFTIN1, SHIFTIN2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input BITSLIP ;
input CE1 ;
input CE2 ;
input CLK ;
input CLKB ;
input CLKDIV ;
input D ;
input DDLY ;
input DYNCLKDIVSEL ;
input DYNCLKSEL ;
input OCLK ;
input OFB ;
input RST ;
input SHIFTIN1 ;
input SHIFTIN2 ;
output O ;
output Q1 ;
output Q2 ;
output Q3 ;
output Q4 ;
output Q5 ;
output Q6 ;
output SHIFTOUT1 ;
output SHIFTOUT2 ;
parameter DATA_RATE = "DDR";
parameter DATA_WIDTH = 4;
parameter DYN_CLKDIV_INV_EN = "FALSE";
parameter DYN_CLK_INV_EN = "FALSE";
parameter INIT_Q1 = 1'b0;
parameter INIT_Q2 = 1'b0;
parameter INIT_Q3 = 1'b0;
parameter INIT_Q4 = 1'b0;
parameter INTERFACE_TYPE = "MEMORY";
parameter NUM_CE = 2;
parameter IOBDELAY = "NONE";
parameter OFB_USED = "FALSE";
parameter SERDES_MODE = "MASTER";
parameter SRVAL_Q1 = 1'b0;
parameter SRVAL_Q2 = 1'b0;
parameter SRVAL_Q3 = 1'b0;
parameter SRVAL_Q4 = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: ISERDESE1 ####

//#### BEGIN MODULE DEFINITION FOR :ISERDESE2 ###
module ISERDESE2 (
  O,
  Q1,
  Q2,
  Q3,
  Q4,
  Q5,
  Q6,
  Q7,
  Q8,
  SHIFTOUT1,
  SHIFTOUT2,

  BITSLIP,
  CE1,
  CE2,
  CLK,
  CLKB,
  CLKDIV,
  CLKDIVP,
  D,
  DDLY,
  DYNCLKDIVSEL,
  DYNCLKSEL,
  OCLK,
  OCLKB,
  OFB,
  RST,
  SHIFTIN1,
  SHIFTIN2
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input BITSLIP ;
input CE1 ;
input CE2 ;
input CLK ;
input CLKB ;
input CLKDIV ;
input CLKDIVP ;
input D ;
input DDLY ;
input DYNCLKDIVSEL ;
input DYNCLKSEL ;
input OCLK ;
input OCLKB ;
input OFB ;
input RST ;
input SHIFTIN1 ;
input SHIFTIN2 ;
output O ;
output Q1 ;
output Q2 ;
output Q3 ;
output Q4 ;
output Q5 ;
output Q6 ;
output Q7 ;
output Q8 ;
output SHIFTOUT1 ;
output SHIFTOUT2 ;
parameter DATA_RATE = "DDR";
parameter DATA_WIDTH = 4;
parameter DYN_CLKDIV_INV_EN = "FALSE";
parameter DYN_CLK_INV_EN = "FALSE";
parameter [0:0] INIT_Q1 = 1'b0;
parameter [0:0] INIT_Q2 = 1'b0;
parameter [0:0] INIT_Q3 = 1'b0;
parameter [0:0] INIT_Q4 = 1'b0;
parameter INTERFACE_TYPE = "MEMORY";
parameter IOBDELAY = "NONE";
parameter NUM_CE = 2;
parameter OFB_USED = "FALSE";
parameter SERDES_MODE = "MASTER";
parameter [0:0] SRVAL_Q1 = 1'b0;
parameter [0:0] SRVAL_Q2 = 1'b0;
parameter [0:0] SRVAL_Q3 = 1'b0;
parameter [0:0] SRVAL_Q4 = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: ISERDESE2 ####

//#### BEGIN MODULE DEFINITION FOR :ISERDES_NODELAY ###
module ISERDES_NODELAY (Q1, Q2, Q3, Q4, Q5, Q6, SHIFTOUT1, SHIFTOUT2,
		  BITSLIP, CE1, CE2, CLK, CLKB, CLKDIV, D, OCLK, RST, SHIFTIN1, SHIFTIN2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input BITSLIP ;
input CE1 ;
input CE2 ;
input CLK ;
input CLKB ;
input CLKDIV ;
input D ;
input OCLK ;
input RST ;
input SHIFTIN1 ;
input SHIFTIN2 ;
output Q1 ;
output Q2 ;
output Q3 ;
output Q4 ;
output Q5 ;
output Q6 ;
output SHIFTOUT1 ;
output SHIFTOUT2 ;
parameter BITSLIP_ENABLE = "FALSE";
parameter DATA_RATE = "DDR";
parameter DATA_WIDTH = 4;
parameter INIT_Q1 = 1'b0;
parameter INIT_Q2 = 1'b0;
parameter INIT_Q3 = 1'b0;
parameter INIT_Q4 = 1'b0;
parameter INTERFACE_TYPE = "MEMORY";
parameter NUM_CE = 2;
parameter SERDES_MODE = "MASTER";
endmodule
//#### END MODULE DEFINITION FOR: ISERDES_NODELAY ####

//#### BEGIN MODULE DEFINITION FOR :JTAGPPC ###
module JTAGPPC (TCK, TDIPPC, TMS, TDOPPC, TDOTSPPC) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input TDOPPC ;
input TDOTSPPC ;
output TCK ;
output TDIPPC ;
output TMS ;
endmodule
//#### END MODULE DEFINITION FOR: JTAGPPC ####

//#### BEGIN MODULE DEFINITION FOR :JTAGPPC440 ###
module JTAGPPC440 (
        TCK,
        TDIPPC,
        TMS,
        TDOPPC
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input TDOPPC ;
output TCK ;
output TDIPPC ;
output TMS ;
endmodule
//#### END MODULE DEFINITION FOR: JTAGPPC440 ####

//#### BEGIN MODULE DEFINITION FOR :JTAG_SIME2 ###
module JTAG_SIME2( TDO, TCK, TDI, TMS) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input TCK ;
input TDI ;
input TMS ;
output TDO ;
parameter PART_NAME = "7A8";
endmodule
//#### END MODULE DEFINITION FOR: JTAG_SIME2 ####

//#### BEGIN MODULE DEFINITION FOR :JTAG_SIM_SPARTAN3A ###
module JTAG_SIM_SPARTAN3A( TDO, TCK, TDI, TMS ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input TCK ;
input TDI ;
input TMS ;
output TDO ;
parameter PART_NAME = "3S200A";
endmodule
//#### END MODULE DEFINITION FOR: JTAG_SIM_SPARTAN3A ####

//#### BEGIN MODULE DEFINITION FOR :JTAG_SIM_SPARTAN6 ###
module JTAG_SIM_SPARTAN6( TDO, TCK, TDI, TMS) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input TCK ;
input TDI ;
input TMS ;
output TDO ;
parameter PART_NAME = "LX4";
endmodule
//#### END MODULE DEFINITION FOR: JTAG_SIM_SPARTAN6 ####

//#### BEGIN MODULE DEFINITION FOR :JTAG_SIM_VIRTEX4 ###
module JTAG_SIM_VIRTEX4( TDO, TCK, TDI, TMS ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input TCK ;
input TDI ;
input TMS ;
output TDO ;
parameter PART_NAME = "LX15";
endmodule
//#### END MODULE DEFINITION FOR: JTAG_SIM_VIRTEX4 ####

//#### BEGIN MODULE DEFINITION FOR :JTAG_SIM_VIRTEX5 ###
module JTAG_SIM_VIRTEX5( TDO, TCK, TDI, TMS ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input TCK ;
input TDI ;
input TMS ;
output TDO ;
parameter PART_NAME = "LX30";
endmodule
//#### END MODULE DEFINITION FOR: JTAG_SIM_VIRTEX5 ####

//#### BEGIN MODULE DEFINITION FOR :JTAG_SIM_VIRTEX6 ###
module JTAG_SIM_VIRTEX6( TDO, TCK, TDI, TMS) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input TCK ;
input TDI ;
input TMS ;
output TDO ;
parameter PART_NAME = "LX75T";
endmodule
//#### END MODULE DEFINITION FOR: JTAG_SIM_VIRTEX6 ####

//#### BEGIN MODULE DEFINITION FOR :KEEPER ###
module KEEPER (O) /* synthesis syn_black_box  syn_lib_cell=1
 .noprune=1
 */;
inout O ;
endmodule
//#### END MODULE DEFINITION FOR: KEEPER ####

//#### BEGIN MODULE DEFINITION FOR :KEY_CLEAR ###
module KEY_CLEAR (
	KEYCLEARB
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input KEYCLEARB ;
endmodule
//#### END MODULE DEFINITION FOR: KEY_CLEAR ####

//#### BEGIN MODULE DEFINITION FOR :LD ###
module LD (Q, D, G) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input D ;
input G ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: LD ####

//#### BEGIN MODULE DEFINITION FOR :LDC ###
module LDC (Q, CLR, D, G) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLR ;
input D ;
input G ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: LDC ####

//#### BEGIN MODULE DEFINITION FOR :LDCE ###
module LDCE (Q, CLR, D, G, GE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLR ;
input D ;
input G ;
input GE ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: LDCE ####

//#### BEGIN MODULE DEFINITION FOR :LDCE_1 ###
module LDCE_1 (Q, CLR, D, G, GE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLR ;
input D ;
input G ;
input GE ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: LDCE_1 ####

//#### BEGIN MODULE DEFINITION FOR :LDCP ###
module LDCP (Q, CLR, D, G, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLR ;
input D ;
input G ;
input PRE ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: LDCP ####

//#### BEGIN MODULE DEFINITION FOR :LDCPE ###
module LDCPE (Q, CLR, D, G, GE, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLR ;
input D ;
input G ;
input GE ;
input PRE ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: LDCPE ####

//#### BEGIN MODULE DEFINITION FOR :LDCPE_1 ###
module LDCPE_1 (Q, CLR, D, G, GE, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLR ;
input D ;
input G ;
input GE ;
input PRE ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: LDCPE_1 ####

//#### BEGIN MODULE DEFINITION FOR :LDCP_1 ###
module LDCP_1 (Q, CLR, D, G, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLR ;
input D ;
input G ;
input PRE ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: LDCP_1 ####

//#### BEGIN MODULE DEFINITION FOR :LDC_1 ###
module LDC_1 (Q, CLR, D, G) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLR ;
input D ;
input G ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: LDC_1 ####

//#### BEGIN MODULE DEFINITION FOR :LDE ###
module LDE (Q, D, G, GE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input D ;
input G ;
input GE ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: LDE ####

//#### BEGIN MODULE DEFINITION FOR :LDE_1 ###
module LDE_1 (Q, D, G, GE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input D ;
input G ;
input GE ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: LDE_1 ####

//#### BEGIN MODULE DEFINITION FOR :LDP ###
module LDP (Q, D, G, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input D ;
input G ;
input PRE ;
output Q ;
parameter INIT = 1'b1;
endmodule
//#### END MODULE DEFINITION FOR: LDP ####

//#### BEGIN MODULE DEFINITION FOR :LDPE ###
module LDPE (Q, D, G, GE, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input D ;
input G ;
input GE ;
input PRE ;
output Q ;
parameter INIT = 1'b1;
endmodule
//#### END MODULE DEFINITION FOR: LDPE ####

//#### BEGIN MODULE DEFINITION FOR :LDPE_1 ###
module LDPE_1 (Q, D, G, GE, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input D ;
input G ;
input GE ;
input PRE ;
output Q ;
parameter INIT = 1'b1;
endmodule
//#### END MODULE DEFINITION FOR: LDPE_1 ####

//#### BEGIN MODULE DEFINITION FOR :LDP_1 ###
module LDP_1 (Q, D, G, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input D ;
input G ;
input PRE ;
output Q ;
parameter INIT = 1'b1;
endmodule
//#### END MODULE DEFINITION FOR: LDP_1 ####

//#### BEGIN MODULE DEFINITION FOR :LD_1 ###
module LD_1 (Q, D, G) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input D ;
input G ;
output Q ;
parameter INIT = 1'b0;
endmodule
//#### END MODULE DEFINITION FOR: LD_1 ####

//#### BEGIN MODULE DEFINITION FOR :LUT1 ###
module LUT1 (O, I0) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
output O ;
parameter INIT = 2'h0;
endmodule
//#### END MODULE DEFINITION FOR: LUT1 ####

//#### BEGIN MODULE DEFINITION FOR :LUT1_D ###
module LUT1_D (LO, O, I0) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
output LO ;
output O ;
parameter INIT = 2'h0;
endmodule
//#### END MODULE DEFINITION FOR: LUT1_D ####

//#### BEGIN MODULE DEFINITION FOR :LUT1_L ###
module LUT1_L (LO, I0) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
output LO ;
parameter INIT = 2'h0;
endmodule
//#### END MODULE DEFINITION FOR: LUT1_L ####

//#### BEGIN MODULE DEFINITION FOR :LUT2 ###
module LUT2 (O, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
input I1 ;
output O ;
parameter INIT = 4'h0;
endmodule
//#### END MODULE DEFINITION FOR: LUT2 ####

//#### BEGIN MODULE DEFINITION FOR :LUT2_D ###
module LUT2_D (LO, O, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
input I1 ;
output LO ;
output O ;
parameter INIT = 4'h0;
endmodule
//#### END MODULE DEFINITION FOR: LUT2_D ####

//#### BEGIN MODULE DEFINITION FOR :LUT2_L ###
module LUT2_L (LO, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
input I1 ;
output LO ;
parameter INIT = 4'h0;
endmodule
//#### END MODULE DEFINITION FOR: LUT2_L ####

//#### BEGIN MODULE DEFINITION FOR :LUT3 ###
module LUT3 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
parameter INIT = 8'h00;
endmodule
//#### END MODULE DEFINITION FOR: LUT3 ####

//#### BEGIN MODULE DEFINITION FOR :LUT3_D ###
module LUT3_D (LO, O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
input I1 ;
input I2 ;
output LO ;
output O ;
parameter INIT = 8'h00;
endmodule
//#### END MODULE DEFINITION FOR: LUT3_D ####

//#### BEGIN MODULE DEFINITION FOR :LUT3_L ###
module LUT3_L (LO, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
input I1 ;
input I2 ;
output LO ;
parameter INIT = 8'h00;
endmodule
//#### END MODULE DEFINITION FOR: LUT3_L ####

//#### BEGIN MODULE DEFINITION FOR :LUT4 ###
module LUT4 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
parameter INIT = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: LUT4 ####

//#### BEGIN MODULE DEFINITION FOR :LUT4_D ###
module LUT4_D (LO, O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
output LO ;
parameter INIT = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: LUT4_D ####

//#### BEGIN MODULE DEFINITION FOR :LUT4_L ###
module LUT4_L (LO, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output LO ;
parameter INIT = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: LUT4_L ####

//#### BEGIN MODULE DEFINITION FOR :LUT5 ###
module LUT5 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
parameter INIT = 32'h00000000;
endmodule
//#### END MODULE DEFINITION FOR: LUT5 ####

//#### BEGIN MODULE DEFINITION FOR :LUT5_D ###
module LUT5_D (LO, O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output LO ;
output O ;
parameter INIT = 32'h00000000;
endmodule
//#### END MODULE DEFINITION FOR: LUT5_D ####

//#### BEGIN MODULE DEFINITION FOR :LUT5_L ###
module LUT5_L (LO, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output LO ;
parameter INIT = 32'h00000000;
endmodule
//#### END MODULE DEFINITION FOR: LUT5_L ####

//#### BEGIN MODULE DEFINITION FOR :LUT6 ###
module LUT6 (O, I0, I1, I2, I3, I4, I5) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
input I5 ;
output O ;
parameter INIT = 64'h0000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: LUT6 ####

//#### BEGIN MODULE DEFINITION FOR :LUT6_2 ###
module LUT6_2 (O5, O6, I0, I1, I2, I3, I4, I5) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
input I5 ;
output O5 ;
output O6 ;
parameter INIT = 64'h0000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: LUT6_2 ####

//#### BEGIN MODULE DEFINITION FOR :LUT6_D ###
module LUT6_D (LO, O, I0, I1, I2, I3, I4, I5) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
input I5 ;
output LO ;
output O ;
parameter INIT = 64'h0000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: LUT6_D ####

//#### BEGIN MODULE DEFINITION FOR :LUT6_L ###
module LUT6_L (LO, I0, I1, I2, I3, I4, I5) /* synthesis syn_black_box  syn_lib_cell=1
 xc_map=lut
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
input I5 ;
output LO ;
parameter INIT = 64'h0000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: LUT6_L ####

//#### BEGIN MODULE DEFINITION FOR :MCB ###
module MCB (
  ADDR,
  BA,
  CAS,
  CKE,
  DQIOWEN0,
  DQON,
  DQOP,
  DQSIOWEN90N,
  DQSIOWEN90P,
  IOIDRPADD,
  IOIDRPADDR,
  IOIDRPBROADCAST,
  IOIDRPCLK,
  IOIDRPCS,
  IOIDRPSDO,
  IOIDRPTRAIN,
  IOIDRPUPDATE,
  LDMN,
  LDMP,
  ODT,
  P0CMDEMPTY,
  P0CMDFULL,
  P0RDCOUNT,
  P0RDDATA,
  P0RDEMPTY,
  P0RDERROR,
  P0RDFULL,
  P0RDOVERFLOW,
  P0WRCOUNT,
  P0WREMPTY,
  P0WRERROR,
  P0WRFULL,
  P0WRUNDERRUN,
  P1CMDEMPTY,
  P1CMDFULL,
  P1RDCOUNT,
  P1RDDATA,
  P1RDEMPTY,
  P1RDERROR,
  P1RDFULL,
  P1RDOVERFLOW,
  P1WRCOUNT,
  P1WREMPTY,
  P1WRERROR,
  P1WRFULL,
  P1WRUNDERRUN,
  P2CMDEMPTY,
  P2CMDFULL,
  P2COUNT,
  P2EMPTY,
  P2ERROR,
  P2FULL,
  P2RDDATA,
  P2RDOVERFLOW,
  P2WRUNDERRUN,
  P3CMDEMPTY,
  P3CMDFULL,
  P3COUNT,
  P3EMPTY,
  P3ERROR,
  P3FULL,
  P3RDDATA,
  P3RDOVERFLOW,
  P3WRUNDERRUN,
  P4CMDEMPTY,
  P4CMDFULL,
  P4COUNT,
  P4EMPTY,
  P4ERROR,
  P4FULL,
  P4RDDATA,
  P4RDOVERFLOW,
  P4WRUNDERRUN,
  P5CMDEMPTY,
  P5CMDFULL,
  P5COUNT,
  P5EMPTY,
  P5ERROR,
  P5FULL,
  P5RDDATA,
  P5RDOVERFLOW,
  P5WRUNDERRUN,
  RAS,
  RST,
  SELFREFRESHMODE,
  STATUS,
  UDMN,
  UDMP,
  UOCALSTART,
  UOCMDREADYIN,
  UODATA,
  UODATAVALID,
  UODONECAL,
  UOREFRSHFLAG,
  UOSDO,
  WE,
  DQI,
  DQSIOIN,
  DQSIOIP,
  IOIDRPSDI,
  P0ARBEN,
  P0CMDBA,
  P0CMDBL,
  P0CMDCA,
  P0CMDCLK,
  P0CMDEN,
  P0CMDINSTR,
  P0CMDRA,
  P0RDCLK,
  P0RDEN,
  P0RWRMASK,
  P0WRCLK,
  P0WRDATA,
  P0WREN,
  P1ARBEN,
  P1CMDBA,
  P1CMDBL,
  P1CMDCA,
  P1CMDCLK,
  P1CMDEN,
  P1CMDINSTR,
  P1CMDRA,
  P1RDCLK,
  P1RDEN,
  P1RWRMASK,
  P1WRCLK,
  P1WRDATA,
  P1WREN,
  P2ARBEN,
  P2CLK,
  P2CMDBA,
  P2CMDBL,
  P2CMDCA,
  P2CMDCLK,
  P2CMDEN,
  P2CMDINSTR,
  P2CMDRA,
  P2EN,
  P2WRDATA,
  P2WRMASK,
  P3ARBEN,
  P3CLK,
  P3CMDBA,
  P3CMDBL,
  P3CMDCA,
  P3CMDCLK,
  P3CMDEN,
  P3CMDINSTR,
  P3CMDRA,
  P3EN,
  P3WRDATA,
  P3WRMASK,
  P4ARBEN,
  P4CLK,
  P4CMDBA,
  P4CMDBL,
  P4CMDCA,
  P4CMDCLK,
  P4CMDEN,
  P4CMDINSTR,
  P4CMDRA,
  P4EN,
  P4WRDATA,
  P4WRMASK,
  P5ARBEN,
  P5CLK,
  P5CMDBA,
  P5CMDBL,
  P5CMDCA,
  P5CMDCLK,
  P5CMDEN,
  P5CMDINSTR,
  P5CMDRA,
  P5EN,
  P5WRDATA,
  P5WRMASK,
  PLLCE,
  PLLCLK,
  PLLLOCK,
  RECAL,
  SELFREFRESHENTER,
  SYSRST,
  UDQSIOIN,
  UDQSIOIP,
  UIADD,
  UIADDR,
  UIBROADCAST,
  UICLK,
  UICMD,
  UICMDEN,
  UICMDIN,
  UICS,
  UIDONECAL,
  UIDQCOUNT,
  UIDQLOWERDEC,
  UIDQLOWERINC,
  UIDQUPPERDEC,
  UIDQUPPERINC,
  UIDRPUPDATE,
  UILDQSDEC,
  UILDQSINC,
  UIREAD,
  UISDI,
  UIUDQSDEC,
  UIUDQSINC
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input DQSIOIN ;
input DQSIOIP ;
input IOIDRPSDI ;
input P0ARBEN ;
input P0CMDCLK ;
input P0CMDEN ;
input P0RDCLK ;
input P0RDEN ;
input P0WRCLK ;
input P0WREN ;
input P1ARBEN ;
input P1CMDCLK ;
input P1CMDEN ;
input P1RDCLK ;
input P1RDEN ;
input P1WRCLK ;
input P1WREN ;
input P2ARBEN ;
input P2CLK ;
input P2CMDCLK ;
input P2CMDEN ;
input P2EN ;
input P3ARBEN ;
input P3CLK ;
input P3CMDCLK ;
input P3CMDEN ;
input P3EN ;
input P4ARBEN ;
input P4CLK ;
input P4CMDCLK ;
input P4CMDEN ;
input P4EN ;
input P5ARBEN ;
input P5CLK ;
input P5CMDCLK ;
input P5CMDEN ;
input P5EN ;
input PLLLOCK ;
input RECAL ;
input SELFREFRESHENTER ;
input SYSRST ;
input UDQSIOIN ;
input UDQSIOIP ;
input UIADD ;
input UIBROADCAST ;
input UICLK ;
input UICMD ;
input UICMDEN ;
input UICMDIN ;
input UICS ;
input UIDONECAL ;
input UIDQLOWERDEC ;
input UIDQLOWERINC ;
input UIDQUPPERDEC ;
input UIDQUPPERINC ;
input UIDRPUPDATE ;
input UILDQSDEC ;
input UILDQSINC ;
input UIREAD ;
input UISDI ;
input UIUDQSDEC ;
input UIUDQSINC ;
input [11:0] P0CMDCA ;
input [11:0] P1CMDCA ;
input [11:0] P2CMDCA ;
input [11:0] P3CMDCA ;
input [11:0] P4CMDCA ;
input [11:0] P5CMDCA ;
input [14:0] P0CMDRA ;
input [14:0] P1CMDRA ;
input [14:0] P2CMDRA ;
input [14:0] P3CMDRA ;
input [14:0] P4CMDRA ;
input [14:0] P5CMDRA ;
input [15:0] DQI ;
input [1:0] PLLCE ;
input [1:0] PLLCLK ;
input [2:0] P0CMDBA ;
input [2:0] P0CMDINSTR ;
input [2:0] P1CMDBA ;
input [2:0] P1CMDINSTR ;
input [2:0] P2CMDBA ;
input [2:0] P2CMDINSTR ;
input [2:0] P3CMDBA ;
input [2:0] P3CMDINSTR ;
input [2:0] P4CMDBA ;
input [2:0] P4CMDINSTR ;
input [2:0] P5CMDBA ;
input [2:0] P5CMDINSTR ;
input [31:0] P0WRDATA ;
input [31:0] P1WRDATA ;
input [31:0] P2WRDATA ;
input [31:0] P3WRDATA ;
input [31:0] P4WRDATA ;
input [31:0] P5WRDATA ;
input [3:0] P0RWRMASK ;
input [3:0] P1RWRMASK ;
input [3:0] P2WRMASK ;
input [3:0] P3WRMASK ;
input [3:0] P4WRMASK ;
input [3:0] P5WRMASK ;
input [3:0] UIDQCOUNT ;
input [4:0] UIADDR ;
input [5:0] P0CMDBL ;
input [5:0] P1CMDBL ;
input [5:0] P2CMDBL ;
input [5:0] P3CMDBL ;
input [5:0] P4CMDBL ;
input [5:0] P5CMDBL ;
output CAS ;
output CKE ;
output DQIOWEN0 ;
output DQSIOWEN90N ;
output DQSIOWEN90P ;
output IOIDRPADD ;
output IOIDRPBROADCAST ;
output IOIDRPCLK ;
output IOIDRPCS ;
output IOIDRPSDO ;
output IOIDRPTRAIN ;
output IOIDRPUPDATE ;
output LDMN ;
output LDMP ;
output ODT ;
output P0CMDEMPTY ;
output P0CMDFULL ;
output P0RDEMPTY ;
output P0RDERROR ;
output P0RDFULL ;
output P0RDOVERFLOW ;
output P0WREMPTY ;
output P0WRERROR ;
output P0WRFULL ;
output P0WRUNDERRUN ;
output P1CMDEMPTY ;
output P1CMDFULL ;
output P1RDEMPTY ;
output P1RDERROR ;
output P1RDFULL ;
output P1RDOVERFLOW ;
output P1WREMPTY ;
output P1WRERROR ;
output P1WRFULL ;
output P1WRUNDERRUN ;
output P2CMDEMPTY ;
output P2CMDFULL ;
output P2EMPTY ;
output P2ERROR ;
output P2FULL ;
output P2RDOVERFLOW ;
output P2WRUNDERRUN ;
output P3CMDEMPTY ;
output P3CMDFULL ;
output P3EMPTY ;
output P3ERROR ;
output P3FULL ;
output P3RDOVERFLOW ;
output P3WRUNDERRUN ;
output P4CMDEMPTY ;
output P4CMDFULL ;
output P4EMPTY ;
output P4ERROR ;
output P4FULL ;
output P4RDOVERFLOW ;
output P4WRUNDERRUN ;
output P5CMDEMPTY ;
output P5CMDFULL ;
output P5EMPTY ;
output P5ERROR ;
output P5FULL ;
output P5RDOVERFLOW ;
output P5WRUNDERRUN ;
output RAS ;
output RST ;
output SELFREFRESHMODE ;
output UDMN ;
output UDMP ;
output UOCALSTART ;
output UOCMDREADYIN ;
output UODATAVALID ;
output UODONECAL ;
output UOREFRSHFLAG ;
output UOSDO ;
output WE ;
output [14:0] ADDR ;
output [15:0] DQON ;
output [15:0] DQOP ;
output [2:0] BA ;
output [31:0] P0RDDATA ;
output [31:0] P1RDDATA ;
output [31:0] P2RDDATA ;
output [31:0] P3RDDATA ;
output [31:0] P4RDDATA ;
output [31:0] P5RDDATA ;
output [31:0] STATUS ;
output [4:0] IOIDRPADDR ;
output [6:0] P0RDCOUNT ;
output [6:0] P0WRCOUNT ;
output [6:0] P1RDCOUNT ;
output [6:0] P1WRCOUNT ;
output [6:0] P2COUNT ;
output [6:0] P3COUNT ;
output [6:0] P4COUNT ;
output [6:0] P5COUNT ;
output [7:0] UODATA ;
parameter ARB_NUM_TIME_SLOTS = 12;
parameter [17:0] ARB_TIME_SLOT_0 = 18'b111111111111111111;
parameter [17:0] ARB_TIME_SLOT_1 = 18'b111111111111111111;
parameter [17:0] ARB_TIME_SLOT_10 = 18'b111111111111111111;
parameter [17:0] ARB_TIME_SLOT_11 = 18'b111111111111111111;
parameter [17:0] ARB_TIME_SLOT_2 = 18'b111111111111111111;
parameter [17:0] ARB_TIME_SLOT_3 = 18'b111111111111111111;
parameter [17:0] ARB_TIME_SLOT_4 = 18'b111111111111111111;
parameter [17:0] ARB_TIME_SLOT_5 = 18'b111111111111111111;
parameter [17:0] ARB_TIME_SLOT_6 = 18'b111111111111111111;
parameter [17:0] ARB_TIME_SLOT_7 = 18'b111111111111111111;
parameter [17:0] ARB_TIME_SLOT_8 = 18'b111111111111111111;
parameter [17:0] ARB_TIME_SLOT_9 = 18'b111111111111111111;
parameter [2:0] CAL_BA = 3'h0;
parameter CAL_BYPASS = "YES";
parameter [11:0] CAL_CA = 12'h000;
parameter CAL_CALIBRATION_MODE = "NOCALIBRATION";
parameter CAL_CLK_DIV = 1;
parameter CAL_DELAY = "QUARTER";
parameter [14:0] CAL_RA = 15'h0000;
parameter MEM_ADDR_ORDER = "BANK_ROW_COLUMN";
parameter MEM_BA_SIZE = 3;
parameter MEM_BURST_LEN = 8;
parameter MEM_CAS_LATENCY = 4;
parameter MEM_CA_SIZE = 11;
parameter MEM_DDR1_2_ODS = "FULL";
parameter MEM_DDR2_3_HIGH_TEMP_SR = "NORMAL";
parameter MEM_DDR2_3_PA_SR = "FULL";
parameter MEM_DDR2_ADD_LATENCY = 0;
parameter MEM_DDR2_DIFF_DQS_EN = "YES";
parameter MEM_DDR2_RTT = "50OHMS";
parameter MEM_DDR2_WRT_RECOVERY = 4;
parameter MEM_DDR3_ADD_LATENCY = "OFF";
parameter MEM_DDR3_AUTO_SR = "ENABLED";
parameter MEM_DDR3_CAS_LATENCY = 7;
parameter MEM_DDR3_CAS_WR_LATENCY = 5;
parameter MEM_DDR3_DYN_WRT_ODT = "OFF";
parameter MEM_DDR3_ODS = "DIV7";
parameter MEM_DDR3_RTT = "DIV2";
parameter MEM_DDR3_WRT_RECOVERY = 7;
parameter MEM_MDDR_ODS = "FULL";
parameter MEM_MOBILE_PA_SR = "FULL";
parameter MEM_MOBILE_TC_SR = 0;
parameter MEM_RAS_VAL = 0;
parameter MEM_RA_SIZE = 13;
parameter MEM_RCD_VAL = 1;
parameter MEM_REFI_VAL = 0;
parameter MEM_RFC_VAL = 0;
parameter MEM_RP_VAL = 0;
parameter MEM_RTP_VAL = 0;
parameter MEM_TYPE = "DDR3";
parameter MEM_WIDTH = 4;
parameter MEM_WR_VAL = 0;
parameter MEM_WTR_VAL = 3;
parameter PORT_CONFIG = "B32_B32_B32_B32";
endmodule
//#### END MODULE DEFINITION FOR: MCB ####

//#### BEGIN MODULE DEFINITION FOR :MMCME2_ADV ###
module MMCME2_ADV (
  CLKFBOUT,
  CLKFBOUTB,
  CLKFBSTOPPED,
  CLKINSTOPPED,
  CLKOUT0,
  CLKOUT0B,
  CLKOUT1,
  CLKOUT1B,
  CLKOUT2,
  CLKOUT2B,
  CLKOUT3,
  CLKOUT3B,
  CLKOUT4,
  CLKOUT5,
  CLKOUT6,
  DO,
  DRDY,
  LOCKED,
  PSDONE,
  CLKFBIN,
  CLKIN1,
  CLKIN2,
  CLKINSEL,
  DADDR,
  DCLK,
  DEN,
  DI,
  DWE,
  PSCLK,
  PSEN,
  PSINCDEC,
  PWRDWN,
  RST
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKFBIN ;
input CLKIN1 ;
input CLKIN2 ;
input CLKINSEL ;
input DCLK ;
input DEN ;
input DWE ;
input PSCLK ;
input PSEN ;
input PSINCDEC ;
input PWRDWN ;
input RST ;
input [15:0] DI ;
input [6:0] DADDR ;
output CLKFBOUT ;
output CLKFBOUTB ;
output CLKFBSTOPPED ;
output CLKINSTOPPED ;
output CLKOUT0 ;
output CLKOUT0B ;
output CLKOUT1 ;
output CLKOUT1B ;
output CLKOUT2 ;
output CLKOUT2B ;
output CLKOUT3 ;
output CLKOUT3B ;
output CLKOUT4 ;
output CLKOUT5 ;
output CLKOUT6 ;
output DRDY ;
output LOCKED ;
output PSDONE ;
output [15:0] DO ;
parameter BANDWIDTH = "OPTIMIZED";
parameter CLKFBOUT_USE_FINE_PS = "FALSE";
parameter CLKOUT0_USE_FINE_PS = "FALSE";
parameter CLKOUT1_USE_FINE_PS = "FALSE";
parameter CLKOUT2_USE_FINE_PS = "FALSE";
parameter CLKOUT3_USE_FINE_PS = "FALSE";
parameter CLKOUT4_CASCADE = "FALSE";
parameter CLKOUT4_USE_FINE_PS = "FALSE";
parameter CLKOUT5_USE_FINE_PS = "FALSE";
parameter CLKOUT6_USE_FINE_PS = "FALSE";
parameter COMPENSATION = "ZHOLD";
parameter STARTUP_WAIT = "FALSE";
parameter CLKOUT1_DIVIDE = 1;
parameter CLKOUT2_DIVIDE = 1;
parameter CLKOUT3_DIVIDE = 1;
parameter CLKOUT4_DIVIDE = 1;
parameter CLKOUT5_DIVIDE = 1;
parameter CLKOUT6_DIVIDE = 1;
parameter DIVCLK_DIVIDE = 1;
parameter CLKFBOUT_MULT_F = 5.000;
parameter CLKFBOUT_PHASE = 0.000;
parameter CLKIN1_PERIOD = 0.000;
parameter CLKIN2_PERIOD = 0.000;
parameter CLKOUT0_DIVIDE_F = 1.000;
parameter CLKOUT0_DUTY_CYCLE = 0.500;
parameter CLKOUT0_PHASE = 0.000;
parameter CLKOUT1_DUTY_CYCLE = 0.500;
parameter CLKOUT1_PHASE = 0.000;
parameter CLKOUT2_DUTY_CYCLE = 0.500;
parameter CLKOUT2_PHASE = 0.000;
parameter CLKOUT3_DUTY_CYCLE = 0.500;
parameter CLKOUT3_PHASE = 0.000;
parameter CLKOUT4_DUTY_CYCLE = 0.500;
parameter CLKOUT4_PHASE = 0.000;
parameter CLKOUT5_DUTY_CYCLE = 0.500;
parameter CLKOUT5_PHASE = 0.000;
parameter CLKOUT6_DUTY_CYCLE = 0.500;
parameter CLKOUT6_PHASE = 0.000;
parameter REF_JITTER1 = 0.010;
parameter REF_JITTER2 = 0.010;
parameter SS_EN = "FALSE";
parameter SS_MODE = "CENTER_HIGH";
parameter SS_MOD_PERIOD = 10000;
endmodule
//#### END MODULE DEFINITION FOR: MMCME2_ADV ####

//#### BEGIN MODULE DEFINITION FOR :MMCME2_BASE ###
module MMCME2_BASE (
  CLKFBOUT,
  CLKFBOUTB,
  CLKOUT0,
  CLKOUT0B,
  CLKOUT1,
  CLKOUT1B,
  CLKOUT2,
  CLKOUT2B,
  CLKOUT3,
  CLKOUT3B,
  CLKOUT4,
  CLKOUT5,
  CLKOUT6,
  LOCKED,
  CLKFBIN,
  CLKIN1,
  PWRDWN,
  RST
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKFBIN ;
input CLKIN1 ;
input PWRDWN ;
input RST ;
output CLKFBOUT ;
output CLKFBOUTB ;
output CLKOUT0 ;
output CLKOUT0B ;
output CLKOUT1 ;
output CLKOUT1B ;
output CLKOUT2 ;
output CLKOUT2B ;
output CLKOUT3 ;
output CLKOUT3B ;
output CLKOUT4 ;
output CLKOUT5 ;
output CLKOUT6 ;
output LOCKED ;
parameter BANDWIDTH = "OPTIMIZED";
parameter CLKFBOUT_MULT_F = 5.000;
parameter CLKFBOUT_PHASE = 0.000;
parameter CLKIN1_PERIOD = 0.000;
parameter CLKOUT0_DIVIDE_F = 1.000;
parameter CLKOUT0_DUTY_CYCLE = 0.500;
parameter CLKOUT0_PHASE = 0.000;
parameter CLKOUT1_DIVIDE = 1;
parameter CLKOUT1_DUTY_CYCLE = 0.500;
parameter CLKOUT1_PHASE = 0.000;
parameter CLKOUT2_DIVIDE = 1;
parameter CLKOUT2_DUTY_CYCLE = 0.500;
parameter CLKOUT2_PHASE = 0.000;
parameter CLKOUT3_DIVIDE = 1;
parameter CLKOUT3_DUTY_CYCLE = 0.500;
parameter CLKOUT3_PHASE = 0.000;
parameter CLKOUT4_CASCADE = "FALSE";
parameter CLKOUT4_DIVIDE = 1;
parameter CLKOUT4_DUTY_CYCLE = 0.500;
parameter CLKOUT4_PHASE = 0.000;
parameter CLKOUT5_DIVIDE = 1;
parameter CLKOUT5_DUTY_CYCLE = 0.500;
parameter CLKOUT5_PHASE = 0.000;
parameter CLKOUT6_DIVIDE = 1;
parameter CLKOUT6_DUTY_CYCLE = 0.500;
parameter CLKOUT6_PHASE = 0.000;
parameter DIVCLK_DIVIDE = 1;
parameter REF_JITTER1 = 0.010;
parameter STARTUP_WAIT = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: MMCME2_BASE ####

//#### BEGIN MODULE DEFINITION FOR :MMCM_ADV ###
module MMCM_ADV (
  CLKFBOUT,
  CLKFBOUTB,
  CLKFBSTOPPED,
  CLKINSTOPPED,
  CLKOUT0,
  CLKOUT0B,
  CLKOUT1,
  CLKOUT1B,
  CLKOUT2,
  CLKOUT2B,
  CLKOUT3,
  CLKOUT3B,
  CLKOUT4,
  CLKOUT5,
  CLKOUT6,
  DO,
  DRDY,
  LOCKED,
  PSDONE,
  CLKFBIN,
  CLKIN1,
  CLKIN2,
  CLKINSEL,
  DADDR,
  DCLK,
  DEN,
  DI,
  DWE,
  PSCLK,
  PSEN,
  PSINCDEC,
  PWRDWN,
  RST
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKFBIN ;
input CLKIN1 ;
input CLKIN2 ;
input CLKINSEL ;
input DCLK ;
input DEN ;
input DWE ;
input PSCLK ;
input PSEN ;
input PSINCDEC ;
input PWRDWN ;
input RST ;
input [15:0] DI ;
input [6:0] DADDR ;
output CLKFBOUT ;
output CLKFBOUTB ;
output CLKFBSTOPPED ;
output CLKINSTOPPED ;
output CLKOUT0 ;
output CLKOUT0B ;
output CLKOUT1 ;
output CLKOUT1B ;
output CLKOUT2 ;
output CLKOUT2B ;
output CLKOUT3 ;
output CLKOUT3B ;
output CLKOUT4 ;
output CLKOUT5 ;
output CLKOUT6 ;
output DRDY ;
output LOCKED ;
output PSDONE ;
output [15:0] DO ;
parameter BANDWIDTH = "OPTIMIZED";
parameter CLKFBOUT_USE_FINE_PS = "FALSE";
parameter CLKOUT0_USE_FINE_PS = "FALSE";
parameter CLKOUT1_USE_FINE_PS = "FALSE";
parameter CLKOUT2_USE_FINE_PS = "FALSE";
parameter CLKOUT3_USE_FINE_PS = "FALSE";
parameter CLKOUT4_CASCADE = "FALSE";
parameter CLKOUT4_USE_FINE_PS = "FALSE";
parameter CLKOUT5_USE_FINE_PS = "FALSE";
parameter CLKOUT6_USE_FINE_PS = "FALSE";
parameter CLOCK_HOLD = "FALSE";
parameter COMPENSATION = "ZHOLD";
parameter STARTUP_WAIT = "FALSE";
parameter CLKOUT1_DIVIDE = 1;
parameter CLKOUT2_DIVIDE = 1;
parameter CLKOUT3_DIVIDE = 1;
parameter CLKOUT4_DIVIDE = 1;
parameter CLKOUT5_DIVIDE = 1;
parameter CLKOUT6_DIVIDE = 1;
parameter DIVCLK_DIVIDE = 1;
parameter CLKFBOUT_MULT_F = 5.000;
parameter CLKFBOUT_PHASE = 0.000;
parameter CLKIN1_PERIOD = 0.000;
parameter CLKIN2_PERIOD = 0.000;
parameter CLKOUT0_DIVIDE_F = 1.000;
parameter CLKOUT0_DUTY_CYCLE = 0.500;
parameter CLKOUT0_PHASE = 0.000;
parameter CLKOUT1_DUTY_CYCLE = 0.500;
parameter CLKOUT1_PHASE = 0.000;
parameter CLKOUT2_DUTY_CYCLE = 0.500;
parameter CLKOUT2_PHASE = 0.000;
parameter CLKOUT3_DUTY_CYCLE = 0.500;
parameter CLKOUT3_PHASE = 0.000;
parameter CLKOUT4_DUTY_CYCLE = 0.500;
parameter CLKOUT4_PHASE = 0.000;
parameter CLKOUT5_DUTY_CYCLE = 0.500;
parameter CLKOUT5_PHASE = 0.000;
parameter CLKOUT6_DUTY_CYCLE = 0.500;
parameter CLKOUT6_PHASE = 0.000;
parameter REF_JITTER1 = 0.010;
parameter REF_JITTER2 = 0.010;
endmodule
//#### END MODULE DEFINITION FOR: MMCM_ADV ####

//#### BEGIN MODULE DEFINITION FOR :MMCM_BASE ###
module MMCM_BASE (
  CLKFBOUT,
  CLKFBOUTB,
  CLKOUT0,
  CLKOUT0B,
  CLKOUT1,
  CLKOUT1B,
  CLKOUT2,
  CLKOUT2B,
  CLKOUT3,
  CLKOUT3B,
  CLKOUT4,
  CLKOUT5,
  CLKOUT6,
  LOCKED,
  CLKFBIN,
  CLKIN1,
  PWRDWN,
  RST
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKFBIN ;
input CLKIN1 ;
input PWRDWN ;
input RST ;
output CLKFBOUT ;
output CLKFBOUTB ;
output CLKOUT0 ;
output CLKOUT0B ;
output CLKOUT1 ;
output CLKOUT1B ;
output CLKOUT2 ;
output CLKOUT2B ;
output CLKOUT3 ;
output CLKOUT3B ;
output CLKOUT4 ;
output CLKOUT5 ;
output CLKOUT6 ;
output LOCKED ;
parameter BANDWIDTH = "OPTIMIZED";
parameter CLKFBOUT_MULT_F = 5.000;
parameter CLKFBOUT_PHASE = 0.000;
parameter CLKIN1_PERIOD = 0.000;
parameter CLKOUT0_DIVIDE_F = 1.000;
parameter CLKOUT0_DUTY_CYCLE = 0.500;
parameter CLKOUT0_PHASE = 0.000;
parameter CLKOUT1_DIVIDE = 1;
parameter CLKOUT1_DUTY_CYCLE = 0.500;
parameter CLKOUT1_PHASE = 0.000;
parameter CLKOUT2_DIVIDE = 1;
parameter CLKOUT2_DUTY_CYCLE = 0.500;
parameter CLKOUT2_PHASE = 0.000;
parameter CLKOUT3_DIVIDE = 1;
parameter CLKOUT3_DUTY_CYCLE = 0.500;
parameter CLKOUT3_PHASE = 0.000;
parameter CLKOUT4_CASCADE = "FALSE";
parameter CLKOUT4_DIVIDE = 1;
parameter CLKOUT4_DUTY_CYCLE = 0.500;
parameter CLKOUT4_PHASE = 0.000;
parameter CLKOUT5_DIVIDE = 1;
parameter CLKOUT5_DUTY_CYCLE = 0.500;
parameter CLKOUT5_PHASE = 0.000;
parameter CLKOUT6_DIVIDE = 1;
parameter CLKOUT6_DUTY_CYCLE = 0.500;
parameter CLKOUT6_PHASE = 0.000;
parameter CLOCK_HOLD = "FALSE";
parameter DIVCLK_DIVIDE = 1;
parameter REF_JITTER1 = 0.010;
parameter STARTUP_WAIT = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: MMCM_BASE ####

//#### BEGIN MODULE DEFINITION FOR :MULT18X18 ###
module MULT18X18 (P, A, B) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [17:0] A ;
input [17:0] B ;
output [35:0] P ;
endmodule
//#### END MODULE DEFINITION FOR: MULT18X18 ####

//#### BEGIN MODULE DEFINITION FOR :MULT18X18S ###
module MULT18X18S (P, A, B, C, CE, R) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [17:0] A ;
input [17:0] B ;
input C ;
input CE ;
input R ;
output [35:0] P ;
endmodule
//#### END MODULE DEFINITION FOR: MULT18X18S ####

//#### BEGIN MODULE DEFINITION FOR :MULT18X18SIO ###
module MULT18X18SIO (BCOUT, P, A, B, BCIN, CEA, CEB, CEP, CLK, RSTA, RSTB, RSTP)  /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [17:0] A ;
input [17:0] B ;
input [17:0] BCIN ;
input CEA ;
input CEB ;
input CEP ;
input CLK ;
input RSTA ;
input RSTB ;
input RSTP ;
output [17:0] BCOUT ;
output [35:0] P ;
parameter AREG = 1;
parameter BREG = 1;
parameter B_INPUT = "DIRECT";
parameter PREG = 1;
endmodule
//#### END MODULE DEFINITION FOR: MULT18X18SIO ####

//#### BEGIN MODULE DEFINITION FOR :MULT_AND ###
module MULT_AND (LO, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
output LO ;
endmodule
//#### END MODULE DEFINITION FOR: MULT_AND ####

//#### BEGIN MODULE DEFINITION FOR :MUXCY ###
module MUXCY (O, CI, DI, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CI ;
input DI ;
input S ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: MUXCY ####

//#### BEGIN MODULE DEFINITION FOR :MUXCY_D ###
module MUXCY_D (LO, O, CI, DI, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CI ;
input DI ;
input S ;
output LO ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: MUXCY_D ####

//#### BEGIN MODULE DEFINITION FOR :MUXCY_L ###
module MUXCY_L (LO, CI, DI, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CI ;
input DI ;
input S ;
output LO ;
endmodule
//#### END MODULE DEFINITION FOR: MUXCY_L ####

//#### BEGIN MODULE DEFINITION FOR :MUXF5 ###
module MUXF5 (O, I0, I1, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input S ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: MUXF5 ####

//#### BEGIN MODULE DEFINITION FOR :MUXF5_D ###
module MUXF5_D (LO, O, I0, I1, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input S ;
output LO ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: MUXF5_D ####

//#### BEGIN MODULE DEFINITION FOR :MUXF5_L ###
module MUXF5_L (LO, I0, I1, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input S ;
output LO ;
endmodule
//#### END MODULE DEFINITION FOR: MUXF5_L ####

//#### BEGIN MODULE DEFINITION FOR :MUXF6 ###
module MUXF6 (O, I0, I1, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input S ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: MUXF6 ####

//#### BEGIN MODULE DEFINITION FOR :MUXF6_D ###
module MUXF6_D (LO, O, I0, I1, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input S ;
output LO ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: MUXF6_D ####

//#### BEGIN MODULE DEFINITION FOR :MUXF6_L ###
module MUXF6_L (LO, I0, I1, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input S ;
output LO ;
endmodule
//#### END MODULE DEFINITION FOR: MUXF6_L ####

//#### BEGIN MODULE DEFINITION FOR :MUXF7 ###
module MUXF7 (O, I0, I1, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input S ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: MUXF7 ####

//#### BEGIN MODULE DEFINITION FOR :MUXF7_D ###
module MUXF7_D (LO, O, I0, I1, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input S ;
output LO ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: MUXF7_D ####

//#### BEGIN MODULE DEFINITION FOR :MUXF7_L ###
module MUXF7_L (LO, I0, I1, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input S ;
output LO ;
endmodule
//#### END MODULE DEFINITION FOR: MUXF7_L ####

//#### BEGIN MODULE DEFINITION FOR :MUXF8 ###
module MUXF8 (O, I0, I1, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input S ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: MUXF8 ####

//#### BEGIN MODULE DEFINITION FOR :MUXF8_D ###
module MUXF8_D (LO, O, I0, I1, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input S ;
output LO ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: MUXF8_D ####

//#### BEGIN MODULE DEFINITION FOR :MUXF8_L ###
module MUXF8_L (LO, I0, I1, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input S ;
output LO ;
endmodule
//#### END MODULE DEFINITION FOR: MUXF8_L ####

//#### BEGIN MODULE DEFINITION FOR :NAND2 ###
module NAND2 (O, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND2 ####

//#### BEGIN MODULE DEFINITION FOR :NAND2B1 ###
module NAND2B1 (O, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND2B1 ####

//#### BEGIN MODULE DEFINITION FOR :NAND2B2 ###
module NAND2B2 (O, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND2B2 ####

//#### BEGIN MODULE DEFINITION FOR :NAND3 ###
module NAND3 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND3 ####

//#### BEGIN MODULE DEFINITION FOR :NAND3B1 ###
module NAND3B1 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND3B1 ####

//#### BEGIN MODULE DEFINITION FOR :NAND3B2 ###
module NAND3B2 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND3B2 ####

//#### BEGIN MODULE DEFINITION FOR :NAND3B3 ###
module NAND3B3 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND3B3 ####

//#### BEGIN MODULE DEFINITION FOR :NAND4 ###
module NAND4 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND4 ####

//#### BEGIN MODULE DEFINITION FOR :NAND4B1 ###
module NAND4B1 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND4B1 ####

//#### BEGIN MODULE DEFINITION FOR :NAND4B2 ###
module NAND4B2 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND4B2 ####

//#### BEGIN MODULE DEFINITION FOR :NAND4B3 ###
module NAND4B3 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND4B3 ####

//#### BEGIN MODULE DEFINITION FOR :NAND4B4 ###
module NAND4B4 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND4B4 ####

//#### BEGIN MODULE DEFINITION FOR :NAND5 ###
module NAND5 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND5 ####

//#### BEGIN MODULE DEFINITION FOR :NAND5B1 ###
module NAND5B1 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND5B1 ####

//#### BEGIN MODULE DEFINITION FOR :NAND5B2 ###
module NAND5B2 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND5B2 ####

//#### BEGIN MODULE DEFINITION FOR :NAND5B3 ###
module NAND5B3 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND5B3 ####

//#### BEGIN MODULE DEFINITION FOR :NAND5B4 ###
module NAND5B4 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND5B4 ####

//#### BEGIN MODULE DEFINITION FOR :NAND5B5 ###
module NAND5B5 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NAND5B5 ####

//#### BEGIN MODULE DEFINITION FOR :NOR2 ###
module NOR2 (O, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR2 ####

//#### BEGIN MODULE DEFINITION FOR :NOR2B1 ###
module NOR2B1 (O, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR2B1 ####

//#### BEGIN MODULE DEFINITION FOR :NOR2B2 ###
module NOR2B2 (O, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR2B2 ####

//#### BEGIN MODULE DEFINITION FOR :NOR3 ###
module NOR3 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR3 ####

//#### BEGIN MODULE DEFINITION FOR :NOR3B1 ###
module NOR3B1 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR3B1 ####

//#### BEGIN MODULE DEFINITION FOR :NOR3B2 ###
module NOR3B2 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR3B2 ####

//#### BEGIN MODULE DEFINITION FOR :NOR3B3 ###
module NOR3B3 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR3B3 ####

//#### BEGIN MODULE DEFINITION FOR :NOR4 ###
module NOR4 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR4 ####

//#### BEGIN MODULE DEFINITION FOR :NOR4B1 ###
module NOR4B1 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR4B1 ####

//#### BEGIN MODULE DEFINITION FOR :NOR4B2 ###
module NOR4B2 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR4B2 ####

//#### BEGIN MODULE DEFINITION FOR :NOR4B3 ###
module NOR4B3 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR4B3 ####

//#### BEGIN MODULE DEFINITION FOR :NOR4B4 ###
module NOR4B4 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR4B4 ####

//#### BEGIN MODULE DEFINITION FOR :NOR5 ###
module NOR5 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR5 ####

//#### BEGIN MODULE DEFINITION FOR :NOR5B1 ###
module NOR5B1 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR5B1 ####

//#### BEGIN MODULE DEFINITION FOR :NOR5B2 ###
module NOR5B2 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR5B2 ####

//#### BEGIN MODULE DEFINITION FOR :NOR5B3 ###
module NOR5B3 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR5B3 ####

//#### BEGIN MODULE DEFINITION FOR :NOR5B4 ###
module NOR5B4 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR5B4 ####

//#### BEGIN MODULE DEFINITION FOR :NOR5B5 ###
module NOR5B5 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: NOR5B5 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF ###
module OBUF (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
parameter CAPACITANCE = "DONT_CARE";
parameter DRIVE = 12;
parameter IOSTANDARD = "DEFAULT";
parameter SLEW = "SLOW";
endmodule
//#### END MODULE DEFINITION FOR: OBUF ####

//#### BEGIN MODULE DEFINITION FOR :OBUFDS ###
module OBUFDS (O, OB, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
output OB ;
parameter CAPACITANCE = "DONT_CARE";
parameter IOSTANDARD = "DEFAULT";
parameter SLEW = "SLOW";
endmodule
//#### END MODULE DEFINITION FOR: OBUFDS ####

//#### BEGIN MODULE DEFINITION FOR :OBUFDS_BLVDS_25 ###
module OBUFDS_BLVDS_25 (O, OB, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
output OB ;
endmodule
//#### END MODULE DEFINITION FOR: OBUFDS_BLVDS_25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFDS_LDT_25 ###
module OBUFDS_LDT_25 (O, OB, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
output OB ;
endmodule
//#### END MODULE DEFINITION FOR: OBUFDS_LDT_25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFDS_LVDSEXT_25 ###
module OBUFDS_LVDSEXT_25 (O, OB, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
output OB ;
endmodule
//#### END MODULE DEFINITION FOR: OBUFDS_LVDSEXT_25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFDS_LVDSEXT_33 ###
module OBUFDS_LVDSEXT_33 (O, OB, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
output OB ;
endmodule
//#### END MODULE DEFINITION FOR: OBUFDS_LVDSEXT_33 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFDS_LVDS_25 ###
module OBUFDS_LVDS_25 (O, OB, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
output OB ;
endmodule
//#### END MODULE DEFINITION FOR: OBUFDS_LVDS_25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFDS_LVDS_33 ###
module OBUFDS_LVDS_33 (O, OB, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
output OB ;
endmodule
//#### END MODULE DEFINITION FOR: OBUFDS_LVDS_33 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFDS_LVPECL_25 ###
module OBUFDS_LVPECL_25 (O, OB, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
output OB ;
endmodule
//#### END MODULE DEFINITION FOR: OBUFDS_LVPECL_25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFDS_LVPECL_33 ###
module OBUFDS_LVPECL_33 (O, OB, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
output OB ;
endmodule
//#### END MODULE DEFINITION FOR: OBUFDS_LVPECL_33 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFDS_ULVDS_25 ###
module OBUFDS_ULVDS_25 (O, OB, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
output OB ;
endmodule
//#### END MODULE DEFINITION FOR: OBUFDS_ULVDS_25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT ###
module OBUFT (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
parameter CAPACITANCE = "DONT_CARE";
parameter DRIVE = 12;
parameter IOSTANDARD = "DEFAULT";
parameter SLEW = "SLOW";
endmodule
//#### END MODULE DEFINITION FOR: OBUFT ####

//#### BEGIN MODULE DEFINITION FOR :OBUFTDS ###
module OBUFTDS (O, OB, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
output OB /*synthesis syn_tristate=1
 */;
parameter CAPACITANCE = "DONT_CARE";
parameter IOSTANDARD = "DEFAULT";
parameter SLEW = "SLOW";
endmodule
//#### END MODULE DEFINITION FOR: OBUFTDS ####

//#### BEGIN MODULE DEFINITION FOR :OBUFTDS_BLVDS_25 ###
module OBUFTDS_BLVDS_25 (O, OB, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
output OB /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFTDS_BLVDS_25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFTDS_LDT_25 ###
module OBUFTDS_LDT_25 (O, OB, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
output OB /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFTDS_LDT_25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFTDS_LVDSEXT_25 ###
module OBUFTDS_LVDSEXT_25 (O, OB, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
output OB /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFTDS_LVDSEXT_25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFTDS_LVDSEXT_33 ###
module OBUFTDS_LVDSEXT_33 (O, OB, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
output OB /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFTDS_LVDSEXT_33 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFTDS_LVDS_25 ###
module OBUFTDS_LVDS_25 (O, OB, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
output OB /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFTDS_LVDS_25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFTDS_LVDS_33 ###
module OBUFTDS_LVDS_33 (O, OB, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
output OB /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFTDS_LVDS_33 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFTDS_LVPECL_25 ###
module OBUFTDS_LVPECL_25 (O, OB, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
output OB /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFTDS_LVPECL_25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFTDS_LVPECL_33 ###
module OBUFTDS_LVPECL_33 (O, OB, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
output OB /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFTDS_LVPECL_33 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFTDS_ULVDS_25 ###
module OBUFTDS_ULVDS_25 (O, OB, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
output OB /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFTDS_ULVDS_25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_AGP ###
module OBUFT_AGP (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_AGP ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_CTT ###
module OBUFT_CTT (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_CTT ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_F_12 ###
module OBUFT_F_12 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_F_16 ###
module OBUFT_F_16 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_F_2 ###
module OBUFT_F_2 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_F_24 ###
module OBUFT_F_24 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_F_24 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_F_4 ###
module OBUFT_F_4 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_F_6 ###
module OBUFT_F_6 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_F_8 ###
module OBUFT_F_8 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_GTL ###
module OBUFT_GTL (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_GTL ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_GTLP ###
module OBUFT_GTLP (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_GTLP ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_GTLP_DCI ###
module OBUFT_GTLP_DCI (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_GTLP_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_GTL_DCI ###
module OBUFT_GTL_DCI (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_GTL_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_HSTL_I ###
module OBUFT_HSTL_I (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_HSTL_I ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_HSTL_II ###
module OBUFT_HSTL_II (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_HSTL_II ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_HSTL_III ###
module OBUFT_HSTL_III (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_HSTL_III ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_HSTL_III_18 ###
module OBUFT_HSTL_III_18 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_HSTL_III_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_HSTL_III_DCI ###
module OBUFT_HSTL_III_DCI (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_HSTL_III_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_HSTL_III_DCI_18 ###
module OBUFT_HSTL_III_DCI_18 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_HSTL_III_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_HSTL_II_18 ###
module OBUFT_HSTL_II_18 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_HSTL_II_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_HSTL_II_DCI ###
module OBUFT_HSTL_II_DCI (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_HSTL_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_HSTL_II_DCI_18 ###
module OBUFT_HSTL_II_DCI_18 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_HSTL_II_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_HSTL_IV ###
module OBUFT_HSTL_IV (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_HSTL_IV ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_HSTL_IV_18 ###
module OBUFT_HSTL_IV_18 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_HSTL_IV_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_HSTL_IV_DCI ###
module OBUFT_HSTL_IV_DCI (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_HSTL_IV_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_HSTL_IV_DCI_18 ###
module OBUFT_HSTL_IV_DCI_18 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_HSTL_IV_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_HSTL_I_18 ###
module OBUFT_HSTL_I_18 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_HSTL_I_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_HSTL_I_DCI ###
module OBUFT_HSTL_I_DCI (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_HSTL_I_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_HSTL_I_DCI_18 ###
module OBUFT_HSTL_I_DCI_18 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_HSTL_I_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS12 ###
module OBUFT_LVCMOS12 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS12_F_2 ###
module OBUFT_LVCMOS12_F_2 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS12_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS12_F_4 ###
module OBUFT_LVCMOS12_F_4 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS12_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS12_F_6 ###
module OBUFT_LVCMOS12_F_6 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS12_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS12_F_8 ###
module OBUFT_LVCMOS12_F_8 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS12_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS12_S_2 ###
module OBUFT_LVCMOS12_S_2 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS12_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS12_S_4 ###
module OBUFT_LVCMOS12_S_4 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS12_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS12_S_6 ###
module OBUFT_LVCMOS12_S_6 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS12_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS12_S_8 ###
module OBUFT_LVCMOS12_S_8 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS12_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS15 ###
module OBUFT_LVCMOS15 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS15 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS15_F_12 ###
module OBUFT_LVCMOS15_F_12 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS15_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS15_F_16 ###
module OBUFT_LVCMOS15_F_16 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS15_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS15_F_2 ###
module OBUFT_LVCMOS15_F_2 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS15_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS15_F_4 ###
module OBUFT_LVCMOS15_F_4 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS15_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS15_F_6 ###
module OBUFT_LVCMOS15_F_6 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS15_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS15_F_8 ###
module OBUFT_LVCMOS15_F_8 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS15_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS15_S_12 ###
module OBUFT_LVCMOS15_S_12 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS15_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS15_S_16 ###
module OBUFT_LVCMOS15_S_16 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS15_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS15_S_2 ###
module OBUFT_LVCMOS15_S_2 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS15_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS15_S_4 ###
module OBUFT_LVCMOS15_S_4 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS15_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS15_S_6 ###
module OBUFT_LVCMOS15_S_6 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS15_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS15_S_8 ###
module OBUFT_LVCMOS15_S_8 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS15_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS18 ###
module OBUFT_LVCMOS18 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS18_F_12 ###
module OBUFT_LVCMOS18_F_12 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS18_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS18_F_16 ###
module OBUFT_LVCMOS18_F_16 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS18_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS18_F_2 ###
module OBUFT_LVCMOS18_F_2 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS18_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS18_F_4 ###
module OBUFT_LVCMOS18_F_4 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS18_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS18_F_6 ###
module OBUFT_LVCMOS18_F_6 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS18_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS18_F_8 ###
module OBUFT_LVCMOS18_F_8 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS18_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS18_S_12 ###
module OBUFT_LVCMOS18_S_12 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS18_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS18_S_16 ###
module OBUFT_LVCMOS18_S_16 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS18_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS18_S_2 ###
module OBUFT_LVCMOS18_S_2 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS18_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS18_S_4 ###
module OBUFT_LVCMOS18_S_4 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS18_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS18_S_6 ###
module OBUFT_LVCMOS18_S_6 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS18_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS18_S_8 ###
module OBUFT_LVCMOS18_S_8 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS18_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS2 ###
module OBUFT_LVCMOS2 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS25 ###
module OBUFT_LVCMOS25 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS25_F_12 ###
module OBUFT_LVCMOS25_F_12 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS25_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS25_F_16 ###
module OBUFT_LVCMOS25_F_16 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS25_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS25_F_2 ###
module OBUFT_LVCMOS25_F_2 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS25_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS25_F_24 ###
module OBUFT_LVCMOS25_F_24 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS25_F_24 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS25_F_4 ###
module OBUFT_LVCMOS25_F_4 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS25_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS25_F_6 ###
module OBUFT_LVCMOS25_F_6 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS25_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS25_F_8 ###
module OBUFT_LVCMOS25_F_8 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS25_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS25_S_12 ###
module OBUFT_LVCMOS25_S_12 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS25_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS25_S_16 ###
module OBUFT_LVCMOS25_S_16 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS25_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS25_S_2 ###
module OBUFT_LVCMOS25_S_2 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS25_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS25_S_24 ###
module OBUFT_LVCMOS25_S_24 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS25_S_24 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS25_S_4 ###
module OBUFT_LVCMOS25_S_4 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS25_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS25_S_6 ###
module OBUFT_LVCMOS25_S_6 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS25_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS25_S_8 ###
module OBUFT_LVCMOS25_S_8 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS25_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS33 ###
module OBUFT_LVCMOS33 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS33 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS33_F_12 ###
module OBUFT_LVCMOS33_F_12 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS33_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS33_F_16 ###
module OBUFT_LVCMOS33_F_16 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS33_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS33_F_2 ###
module OBUFT_LVCMOS33_F_2 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS33_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS33_F_24 ###
module OBUFT_LVCMOS33_F_24 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS33_F_24 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS33_F_4 ###
module OBUFT_LVCMOS33_F_4 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS33_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS33_F_6 ###
module OBUFT_LVCMOS33_F_6 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS33_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS33_F_8 ###
module OBUFT_LVCMOS33_F_8 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS33_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS33_S_12 ###
module OBUFT_LVCMOS33_S_12 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS33_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS33_S_16 ###
module OBUFT_LVCMOS33_S_16 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS33_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS33_S_2 ###
module OBUFT_LVCMOS33_S_2 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS33_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS33_S_24 ###
module OBUFT_LVCMOS33_S_24 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS33_S_24 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS33_S_4 ###
module OBUFT_LVCMOS33_S_4 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS33_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS33_S_6 ###
module OBUFT_LVCMOS33_S_6 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS33_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVCMOS33_S_8 ###
module OBUFT_LVCMOS33_S_8 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVCMOS33_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVDCI_15 ###
module OBUFT_LVDCI_15 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVDCI_15 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVDCI_18 ###
module OBUFT_LVDCI_18 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVDCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVDCI_25 ###
module OBUFT_LVDCI_25 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVDCI_25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVDCI_33 ###
module OBUFT_LVDCI_33 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVDCI_33 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVDCI_DV2_15 ###
module OBUFT_LVDCI_DV2_15 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVDCI_DV2_15 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVDCI_DV2_18 ###
module OBUFT_LVDCI_DV2_18 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVDCI_DV2_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVDCI_DV2_25 ###
module OBUFT_LVDCI_DV2_25 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVDCI_DV2_25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVDCI_DV2_33 ###
module OBUFT_LVDCI_DV2_33 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVDCI_DV2_33 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVDS ###
module OBUFT_LVDS (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVDS ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVPECL ###
module OBUFT_LVPECL (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVPECL ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVTTL ###
module OBUFT_LVTTL (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVTTL ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVTTL_F_12 ###
module OBUFT_LVTTL_F_12 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVTTL_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVTTL_F_16 ###
module OBUFT_LVTTL_F_16 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVTTL_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVTTL_F_2 ###
module OBUFT_LVTTL_F_2 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVTTL_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVTTL_F_24 ###
module OBUFT_LVTTL_F_24 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVTTL_F_24 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVTTL_F_4 ###
module OBUFT_LVTTL_F_4 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVTTL_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVTTL_F_6 ###
module OBUFT_LVTTL_F_6 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVTTL_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVTTL_F_8 ###
module OBUFT_LVTTL_F_8 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVTTL_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVTTL_S_12 ###
module OBUFT_LVTTL_S_12 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVTTL_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVTTL_S_16 ###
module OBUFT_LVTTL_S_16 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVTTL_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVTTL_S_2 ###
module OBUFT_LVTTL_S_2 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVTTL_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVTTL_S_24 ###
module OBUFT_LVTTL_S_24 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVTTL_S_24 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVTTL_S_4 ###
module OBUFT_LVTTL_S_4 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVTTL_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVTTL_S_6 ###
module OBUFT_LVTTL_S_6 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVTTL_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_LVTTL_S_8 ###
module OBUFT_LVTTL_S_8 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_LVTTL_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_PCI33_3 ###
module OBUFT_PCI33_3 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_PCI33_3 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_PCI33_5 ###
module OBUFT_PCI33_5 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_PCI33_5 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_PCI66_3 ###
module OBUFT_PCI66_3 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_PCI66_3 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_PCIX ###
module OBUFT_PCIX (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_PCIX ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_PCIX66_3 ###
module OBUFT_PCIX66_3 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_PCIX66_3 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_SSTL18_I ###
module OBUFT_SSTL18_I (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_SSTL18_I ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_SSTL18_II ###
module OBUFT_SSTL18_II (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_SSTL18_II ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_SSTL18_II_DCI ###
module OBUFT_SSTL18_II_DCI (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_SSTL18_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_SSTL18_I_DCI ###
module OBUFT_SSTL18_I_DCI (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_SSTL18_I_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_SSTL2_I ###
module OBUFT_SSTL2_I (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_SSTL2_I ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_SSTL2_II ###
module OBUFT_SSTL2_II (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_SSTL2_II ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_SSTL2_II_DCI ###
module OBUFT_SSTL2_II_DCI (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_SSTL2_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_SSTL2_I_DCI ###
module OBUFT_SSTL2_I_DCI (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_SSTL2_I_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_SSTL3_I ###
module OBUFT_SSTL3_I (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_SSTL3_I ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_SSTL3_II ###
module OBUFT_SSTL3_II (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_SSTL3_II ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_SSTL3_II_DCI ###
module OBUFT_SSTL3_II_DCI (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_SSTL3_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_SSTL3_I_DCI ###
module OBUFT_SSTL3_I_DCI (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_SSTL3_I_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_S_12 ###
module OBUFT_S_12 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_S_16 ###
module OBUFT_S_16 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_S_2 ###
module OBUFT_S_2 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_S_24 ###
module OBUFT_S_24 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_S_24 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_S_4 ###
module OBUFT_S_4 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_S_6 ###
module OBUFT_S_6 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUFT_S_8 ###
module OBUFT_S_8 (O, I, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
input T ;
output O /*synthesis syn_tristate=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: OBUFT_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_AGP ###
module OBUF_AGP (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_AGP ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_CTT ###
module OBUF_CTT (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_CTT ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_F_12 ###
module OBUF_F_12 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_F_16 ###
module OBUF_F_16 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_F_2 ###
module OBUF_F_2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_F_24 ###
module OBUF_F_24 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_F_24 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_F_4 ###
module OBUF_F_4 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_F_6 ###
module OBUF_F_6 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_F_8 ###
module OBUF_F_8 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_GTL ###
module OBUF_GTL (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_GTL ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_GTLP ###
module OBUF_GTLP (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_GTLP ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_GTLP_DCI ###
module OBUF_GTLP_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_GTLP_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_GTL_DCI ###
module OBUF_GTL_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_GTL_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_HSTL_I ###
module OBUF_HSTL_I (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_HSTL_I ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_HSTL_II ###
module OBUF_HSTL_II (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_HSTL_II ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_HSTL_III ###
module OBUF_HSTL_III (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_HSTL_III ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_HSTL_III_18 ###
module OBUF_HSTL_III_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_HSTL_III_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_HSTL_III_DCI ###
module OBUF_HSTL_III_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_HSTL_III_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_HSTL_III_DCI_18 ###
module OBUF_HSTL_III_DCI_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_HSTL_III_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_HSTL_II_18 ###
module OBUF_HSTL_II_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_HSTL_II_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_HSTL_II_DCI ###
module OBUF_HSTL_II_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_HSTL_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_HSTL_II_DCI_18 ###
module OBUF_HSTL_II_DCI_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_HSTL_II_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_HSTL_IV ###
module OBUF_HSTL_IV (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_HSTL_IV ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_HSTL_IV_18 ###
module OBUF_HSTL_IV_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_HSTL_IV_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_HSTL_IV_DCI ###
module OBUF_HSTL_IV_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_HSTL_IV_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_HSTL_IV_DCI_18 ###
module OBUF_HSTL_IV_DCI_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_HSTL_IV_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_HSTL_I_18 ###
module OBUF_HSTL_I_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_HSTL_I_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_HSTL_I_DCI ###
module OBUF_HSTL_I_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_HSTL_I_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_HSTL_I_DCI_18 ###
module OBUF_HSTL_I_DCI_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_HSTL_I_DCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS12 ###
module OBUF_LVCMOS12 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS12_F_2 ###
module OBUF_LVCMOS12_F_2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS12_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS12_F_4 ###
module OBUF_LVCMOS12_F_4 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS12_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS12_F_6 ###
module OBUF_LVCMOS12_F_6 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS12_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS12_F_8 ###
module OBUF_LVCMOS12_F_8 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS12_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS12_S_2 ###
module OBUF_LVCMOS12_S_2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS12_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS12_S_4 ###
module OBUF_LVCMOS12_S_4 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS12_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS12_S_6 ###
module OBUF_LVCMOS12_S_6 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS12_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS12_S_8 ###
module OBUF_LVCMOS12_S_8 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS12_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS15 ###
module OBUF_LVCMOS15 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS15 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS15_F_12 ###
module OBUF_LVCMOS15_F_12 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS15_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS15_F_16 ###
module OBUF_LVCMOS15_F_16 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS15_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS15_F_2 ###
module OBUF_LVCMOS15_F_2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS15_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS15_F_4 ###
module OBUF_LVCMOS15_F_4 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS15_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS15_F_6 ###
module OBUF_LVCMOS15_F_6 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS15_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS15_F_8 ###
module OBUF_LVCMOS15_F_8 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS15_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS15_S_12 ###
module OBUF_LVCMOS15_S_12 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS15_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS15_S_16 ###
module OBUF_LVCMOS15_S_16 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS15_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS15_S_2 ###
module OBUF_LVCMOS15_S_2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS15_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS15_S_4 ###
module OBUF_LVCMOS15_S_4 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS15_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS15_S_6 ###
module OBUF_LVCMOS15_S_6 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS15_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS15_S_8 ###
module OBUF_LVCMOS15_S_8 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS15_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS18 ###
module OBUF_LVCMOS18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS18_F_12 ###
module OBUF_LVCMOS18_F_12 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS18_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS18_F_16 ###
module OBUF_LVCMOS18_F_16 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS18_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS18_F_2 ###
module OBUF_LVCMOS18_F_2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS18_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS18_F_4 ###
module OBUF_LVCMOS18_F_4 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS18_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS18_F_6 ###
module OBUF_LVCMOS18_F_6 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS18_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS18_F_8 ###
module OBUF_LVCMOS18_F_8 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS18_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS18_S_12 ###
module OBUF_LVCMOS18_S_12 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS18_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS18_S_16 ###
module OBUF_LVCMOS18_S_16 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS18_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS18_S_2 ###
module OBUF_LVCMOS18_S_2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS18_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS18_S_4 ###
module OBUF_LVCMOS18_S_4 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS18_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS18_S_6 ###
module OBUF_LVCMOS18_S_6 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS18_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS18_S_8 ###
module OBUF_LVCMOS18_S_8 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS18_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS2 ###
module OBUF_LVCMOS2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS25 ###
module OBUF_LVCMOS25 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS25_F_12 ###
module OBUF_LVCMOS25_F_12 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS25_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS25_F_16 ###
module OBUF_LVCMOS25_F_16 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS25_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS25_F_2 ###
module OBUF_LVCMOS25_F_2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS25_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS25_F_24 ###
module OBUF_LVCMOS25_F_24 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS25_F_24 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS25_F_4 ###
module OBUF_LVCMOS25_F_4 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS25_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS25_F_6 ###
module OBUF_LVCMOS25_F_6 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS25_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS25_F_8 ###
module OBUF_LVCMOS25_F_8 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS25_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS25_S_12 ###
module OBUF_LVCMOS25_S_12 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS25_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS25_S_16 ###
module OBUF_LVCMOS25_S_16 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS25_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS25_S_2 ###
module OBUF_LVCMOS25_S_2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS25_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS25_S_24 ###
module OBUF_LVCMOS25_S_24 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS25_S_24 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS25_S_4 ###
module OBUF_LVCMOS25_S_4 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS25_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS25_S_6 ###
module OBUF_LVCMOS25_S_6 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS25_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS25_S_8 ###
module OBUF_LVCMOS25_S_8 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS25_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS33 ###
module OBUF_LVCMOS33 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS33 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS33_F_12 ###
module OBUF_LVCMOS33_F_12 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS33_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS33_F_16 ###
module OBUF_LVCMOS33_F_16 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS33_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS33_F_2 ###
module OBUF_LVCMOS33_F_2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS33_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS33_F_24 ###
module OBUF_LVCMOS33_F_24 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS33_F_24 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS33_F_4 ###
module OBUF_LVCMOS33_F_4 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS33_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS33_F_6 ###
module OBUF_LVCMOS33_F_6 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS33_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS33_F_8 ###
module OBUF_LVCMOS33_F_8 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS33_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS33_S_12 ###
module OBUF_LVCMOS33_S_12 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS33_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS33_S_16 ###
module OBUF_LVCMOS33_S_16 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS33_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS33_S_2 ###
module OBUF_LVCMOS33_S_2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS33_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS33_S_24 ###
module OBUF_LVCMOS33_S_24 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS33_S_24 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS33_S_4 ###
module OBUF_LVCMOS33_S_4 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS33_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS33_S_6 ###
module OBUF_LVCMOS33_S_6 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS33_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVCMOS33_S_8 ###
module OBUF_LVCMOS33_S_8 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVCMOS33_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVDCI_15 ###
module OBUF_LVDCI_15 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVDCI_15 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVDCI_18 ###
module OBUF_LVDCI_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVDCI_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVDCI_25 ###
module OBUF_LVDCI_25 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVDCI_25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVDCI_33 ###
module OBUF_LVDCI_33 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVDCI_33 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVDCI_DV2_15 ###
module OBUF_LVDCI_DV2_15 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVDCI_DV2_15 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVDCI_DV2_18 ###
module OBUF_LVDCI_DV2_18 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVDCI_DV2_18 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVDCI_DV2_25 ###
module OBUF_LVDCI_DV2_25 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVDCI_DV2_25 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVDCI_DV2_33 ###
module OBUF_LVDCI_DV2_33 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVDCI_DV2_33 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVDS ###
module OBUF_LVDS (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVDS ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVPECL ###
module OBUF_LVPECL (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVPECL ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVTTL ###
module OBUF_LVTTL (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVTTL ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVTTL_F_12 ###
module OBUF_LVTTL_F_12 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVTTL_F_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVTTL_F_16 ###
module OBUF_LVTTL_F_16 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVTTL_F_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVTTL_F_2 ###
module OBUF_LVTTL_F_2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVTTL_F_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVTTL_F_24 ###
module OBUF_LVTTL_F_24 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVTTL_F_24 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVTTL_F_4 ###
module OBUF_LVTTL_F_4 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVTTL_F_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVTTL_F_6 ###
module OBUF_LVTTL_F_6 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVTTL_F_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVTTL_F_8 ###
module OBUF_LVTTL_F_8 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVTTL_F_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVTTL_S_12 ###
module OBUF_LVTTL_S_12 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVTTL_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVTTL_S_16 ###
module OBUF_LVTTL_S_16 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVTTL_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVTTL_S_2 ###
module OBUF_LVTTL_S_2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVTTL_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVTTL_S_24 ###
module OBUF_LVTTL_S_24 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVTTL_S_24 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVTTL_S_4 ###
module OBUF_LVTTL_S_4 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVTTL_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVTTL_S_6 ###
module OBUF_LVTTL_S_6 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVTTL_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_LVTTL_S_8 ###
module OBUF_LVTTL_S_8 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_LVTTL_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_PCI33_3 ###
module OBUF_PCI33_3 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_PCI33_3 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_PCI33_5 ###
module OBUF_PCI33_5 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_PCI33_5 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_PCI66_3 ###
module OBUF_PCI66_3 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_PCI66_3 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_PCIX ###
module OBUF_PCIX (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_PCIX ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_PCIX66_3 ###
module OBUF_PCIX66_3 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_PCIX66_3 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_SSTL18_I ###
module OBUF_SSTL18_I (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_SSTL18_I ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_SSTL18_II ###
module OBUF_SSTL18_II (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_SSTL18_II ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_SSTL18_II_DCI ###
module OBUF_SSTL18_II_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_SSTL18_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_SSTL18_I_DCI ###
module OBUF_SSTL18_I_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_SSTL18_I_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_SSTL2_I ###
module OBUF_SSTL2_I (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_SSTL2_I ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_SSTL2_II ###
module OBUF_SSTL2_II (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_SSTL2_II ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_SSTL2_II_DCI ###
module OBUF_SSTL2_II_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_SSTL2_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_SSTL2_I_DCI ###
module OBUF_SSTL2_I_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_SSTL2_I_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_SSTL3_I ###
module OBUF_SSTL3_I (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_SSTL3_I ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_SSTL3_II ###
module OBUF_SSTL3_II (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_SSTL3_II ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_SSTL3_II_DCI ###
module OBUF_SSTL3_II_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_SSTL3_II_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_SSTL3_I_DCI ###
module OBUF_SSTL3_I_DCI (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_SSTL3_I_DCI ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_S_12 ###
module OBUF_S_12 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_S_12 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_S_16 ###
module OBUF_S_16 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_S_16 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_S_2 ###
module OBUF_S_2 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_S_2 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_S_24 ###
module OBUF_S_24 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_S_24 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_S_4 ###
module OBUF_S_4 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_S_4 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_S_6 ###
module OBUF_S_6 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_S_6 ####

//#### BEGIN MODULE DEFINITION FOR :OBUF_S_8 ###
module OBUF_S_8 (O, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OBUF_S_8 ####

//#### BEGIN MODULE DEFINITION FOR :ODDR ###
module ODDR (Q, C, CE, D1, D2, R, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input D1 ;
input D2 ;
input R ;
input S ;
output Q ;
parameter DDR_CLK_EDGE = "OPPOSITE_EDGE";
parameter INIT = 1'b0;
parameter SRTYPE = "SYNC";
endmodule
//#### END MODULE DEFINITION FOR: ODDR ####

//#### BEGIN MODULE DEFINITION FOR :ODDR2 ###
module ODDR2 (Q, C0, C1, CE, D0, D1, R, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C0 ;
input C1 ;
input CE ;
input D0 ;
input D1 ;
input R ;
input S ;
output Q ;
parameter DDR_ALIGNMENT = "NONE";
parameter INIT = 1'b0;
parameter SRTYPE = "SYNC";
endmodule
//#### END MODULE DEFINITION FOR: ODDR2 ####

//#### BEGIN MODULE DEFINITION FOR :ODELAYE2 ###
module ODELAYE2 (CNTVALUEOUT, DATAOUT, C, CE, CINVCTRL, CLKIN, CNTVALUEIN, INC, LD, LDPIPEEN, ODATAIN, REGRST) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input CINVCTRL ;
input CLKIN ;
input [4:0] CNTVALUEIN ;
input INC ;
input LD ;
input LDPIPEEN ;
input ODATAIN ;
input REGRST ;
output [4:0] CNTVALUEOUT ;
output DATAOUT ;
parameter CINVCTRL_SEL = "FALSE";
parameter DELAY_SRC = "ODATAIN";
parameter HIGH_PERFORMANCE_MODE    = "FALSE";
parameter ODELAY_TYPE  = "FIXED";
parameter ODELAY_VALUE = 0;
parameter PIPE_SEL = "FALSE";
parameter REFCLK_FREQUENCY = 200.0;
parameter SIGNAL_PATTERN    = "DATA";
endmodule
//#### END MODULE DEFINITION FOR: ODELAYE2 ####

//#### BEGIN MODULE DEFINITION FOR :ODELAYE2_FINEDELAY ###
module ODELAYE2_FINEDELAY (
  CNTVALUEOUT,
  DATAOUT,

  C,
  CE,
  CINVCTRL,
  CLKIN,
  CNTVALUEIN,
  INC,
  LD,
  LDPIPEEN,
  ODATAIN,
  OFDLY,
  REGRST
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C ;
input CE ;
input CINVCTRL ;
input CLKIN ;
input [4:0] CNTVALUEIN ;
input INC ;
input LD ;
input LDPIPEEN ;
input ODATAIN ;
input [2:0] OFDLY ;
input REGRST ;
output [4:0] CNTVALUEOUT ;
output DATAOUT ;
parameter CINVCTRL_SEL = "FALSE";
parameter DELAY_SRC = "ODATAIN";
parameter FINEDELAY = "BYPASS";
parameter HIGH_PERFORMANCE_MODE    = "FALSE";
parameter ODELAY_TYPE  = "FIXED";
parameter ODELAY_VALUE = 0;
parameter PIPE_SEL = "FALSE";
parameter REFCLK_FREQUENCY = 200.0;
parameter SIGNAL_PATTERN    = "DATA";
endmodule
//#### END MODULE DEFINITION FOR: ODELAYE2_FINEDELAY ####

//#### BEGIN MODULE DEFINITION FOR :OFDDRCPE ###
module OFDDRCPE (Q, C0, C1, CE, CLR, D0, D1, PRE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C0 ;
input C1 ;
input CE ;
input CLR ;
input D0 ;
input D1 ;
input PRE ;
output Q ;
endmodule
//#### END MODULE DEFINITION FOR: OFDDRCPE ####

//#### BEGIN MODULE DEFINITION FOR :OFDDRRSE ###
module OFDDRRSE (Q, C0, C1, CE, D0, D1, R, S) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C0 ;
input C1 ;
input CE ;
input D0 ;
input D1 ;
input R ;
input S ;
output Q ;
endmodule
//#### END MODULE DEFINITION FOR: OFDDRRSE ####

//#### BEGIN MODULE DEFINITION FOR :OFDDRTCPE ###
module OFDDRTCPE (O, C0, C1, CE, CLR, D0, D1, PRE, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C0 ;
input C1 ;
input CE ;
input CLR ;
input D0 ;
input D1 ;
input PRE ;
input T ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OFDDRTCPE ####

//#### BEGIN MODULE DEFINITION FOR :OFDDRTRSE ###
module OFDDRTRSE (O, C0, C1, CE, D0, D1, R, S, T) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input C0 ;
input C1 ;
input CE ;
input D0 ;
input D1 ;
input R ;
input S ;
input T ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OFDDRTRSE ####

//#### BEGIN MODULE DEFINITION FOR :OR2 ###
module OR2 (O, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR2 ####

//#### BEGIN MODULE DEFINITION FOR :OR2B1 ###
module OR2B1 (O, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR2B1 ####

//#### BEGIN MODULE DEFINITION FOR :OR2B2 ###
module OR2B2 (O, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR2B2 ####

//#### BEGIN MODULE DEFINITION FOR :OR2L ###
module OR2L (O, DI, SRI) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input SRI ;
input DI ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR2L ####

//#### BEGIN MODULE DEFINITION FOR :OR3 ###
module OR3 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR3 ####

//#### BEGIN MODULE DEFINITION FOR :OR3B1 ###
module OR3B1 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR3B1 ####

//#### BEGIN MODULE DEFINITION FOR :OR3B2 ###
module OR3B2 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR3B2 ####

//#### BEGIN MODULE DEFINITION FOR :OR3B3 ###
module OR3B3 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR3B3 ####

//#### BEGIN MODULE DEFINITION FOR :OR4 ###
module OR4 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR4 ####

//#### BEGIN MODULE DEFINITION FOR :OR4B1 ###
module OR4B1 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR4B1 ####

//#### BEGIN MODULE DEFINITION FOR :OR4B2 ###
module OR4B2 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR4B2 ####

//#### BEGIN MODULE DEFINITION FOR :OR4B3 ###
module OR4B3 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR4B3 ####

//#### BEGIN MODULE DEFINITION FOR :OR4B4 ###
module OR4B4 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR4B4 ####

//#### BEGIN MODULE DEFINITION FOR :OR5 ###
module OR5 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR5 ####

//#### BEGIN MODULE DEFINITION FOR :OR5B1 ###
module OR5B1 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR5B1 ####

//#### BEGIN MODULE DEFINITION FOR :OR5B2 ###
module OR5B2 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR5B2 ####

//#### BEGIN MODULE DEFINITION FOR :OR5B3 ###
module OR5B3 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR5B3 ####

//#### BEGIN MODULE DEFINITION FOR :OR5B4 ###
module OR5B4 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR5B4 ####

//#### BEGIN MODULE DEFINITION FOR :OR5B5 ###
module OR5B5 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: OR5B5 ####

//#### BEGIN MODULE DEFINITION FOR :ORCY ###
module ORCY (O, CI, I) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CI ;
input I ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: ORCY ####

//#### BEGIN MODULE DEFINITION FOR :OSERDES ###
module OSERDES (OQ, SHIFTOUT1, SHIFTOUT2, TQ,
		  CLK, CLKDIV, D1, D2, D3, D4, D5, D6, OCE, REV, SHIFTIN1, SHIFTIN2, SR, T1, T2, T3, T4, TCE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLK ;
input CLKDIV ;
input D1 ;
input D2 ;
input D3 ;
input D4 ;
input D5 ;
input D6 ;
input OCE ;
input REV ;
input SHIFTIN1 ;
input SHIFTIN2 ;
input SR ;
input T1 ;
input T2 ;
input T3 ;
input T4 ;
input TCE ;
output OQ ;
output SHIFTOUT1 ;
output SHIFTOUT2 ;
output TQ ;
parameter DATA_RATE_OQ = "DDR";
parameter DATA_RATE_TQ = "DDR";
parameter DATA_WIDTH = 4;
parameter INIT_OQ = 1'b0;
parameter INIT_TQ = 1'b0;
parameter SERDES_MODE = "MASTER";
parameter SRVAL_OQ = 1'b0;
parameter SRVAL_TQ = 1'b0;
parameter TRISTATE_WIDTH = 4;
endmodule
//#### END MODULE DEFINITION FOR: OSERDES ####

//#### BEGIN MODULE DEFINITION FOR :OSERDES2 ###
module OSERDES2 (
  OQ,
  SHIFTOUT1,
  SHIFTOUT2,
  SHIFTOUT3,
  SHIFTOUT4,
  TQ,
  CLK0,
  CLK1,
  CLKDIV,
  D1,
  D2,
  D3,
  D4,
  IOCE,
  OCE,
  RST,
  SHIFTIN1,
  SHIFTIN2,
  SHIFTIN3,
  SHIFTIN4,
  T1,
  T2,
  T3,
  T4,
  TCE,
  TRAIN
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLK0 ;
input CLK1 ;
input CLKDIV ;
input D1 ;
input D2 ;
input D3 ;
input D4 ;
input IOCE ;
input OCE ;
input RST ;
input SHIFTIN1 ;
input SHIFTIN2 ;
input SHIFTIN3 ;
input SHIFTIN4 ;
input T1 ;
input T2 ;
input T3 ;
input T4 ;
input TCE ;
input TRAIN ;
output OQ ;
output SHIFTOUT1 ;
output SHIFTOUT2 ;
output SHIFTOUT3 ;
output SHIFTOUT4 ;
output TQ ;
//output _mode_err_flag= 1 ;
parameter BYPASS_GCLK_FF = "FALSE";
parameter DATA_RATE_OQ = "DDR";
parameter DATA_RATE_OT = "DDR";
parameter DATA_WIDTH =   2;
parameter OUTPUT_MODE = "SINGLE_ENDED";
parameter SERDES_MODE = "NONE";
parameter TRAIN_PATTERN =  0;
endmodule
//#### END MODULE DEFINITION FOR: OSERDES2 ####

//#### BEGIN MODULE DEFINITION FOR :OSERDESE1 ###
module OSERDESE1 (OCBEXTEND, OFB, OQ, SHIFTOUT1, SHIFTOUT2, TFB, TQ,
                    CLK, CLKDIV, CLKPERF, CLKPERFDELAY, D1, D2, D3, D4, D5, D6, OCE, ODV, RST, SHIFTIN1, SHIFTIN2, T1, T2, T3, T4, TCE, WC) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLK ;
input CLKDIV ;
input CLKPERF ;
input CLKPERFDELAY ;
input D1 ;
input D2 ;
input D3 ;
input D4 ;
input D5 ;
input D6 ;
input OCE ;
input ODV ;
input RST ;
input SHIFTIN1 ;
input SHIFTIN2 ;
input T1 ;
input T2 ;
input T3 ;
input T4 ;
input TCE ;
input WC ;
output OCBEXTEND ;
output OFB ;
output OQ ;
output SHIFTOUT1 ;
output SHIFTOUT2 ;
output TFB ;
output TQ ;
parameter DATA_RATE_OQ = "DDR";
parameter DATA_RATE_TQ = "DDR";
parameter DATA_WIDTH = 4;
parameter DDR3_DATA = 1;
parameter INIT_OQ = 1'b0;
parameter INIT_TQ = 1'b0;
parameter INTERFACE_TYPE = "DEFAULT";
parameter ODELAY_USED = 0;
parameter SERDES_MODE = "MASTER";
parameter SRVAL_OQ = 1'b0;
parameter SRVAL_TQ = 1'b0;
parameter TRISTATE_WIDTH = 4;
endmodule
//#### END MODULE DEFINITION FOR: OSERDESE1 ####

//#### BEGIN MODULE DEFINITION FOR :OSERDESE2 ###
module OSERDESE2 (
  OFB,
  OQ,
  SHIFTOUT1,
  SHIFTOUT2,
  TBYTEOUT,
  TFB,
  TQ,

  CLK,
  CLKDIV,
  D1,
  D2,
  D3,
  D4,
  D5,
  D6,
  D7,
  D8,
  OCE,
  RST,
  SHIFTIN1,
  SHIFTIN2,
  T1,
  T2,
  T3,
  T4,
  TBYTEIN,
  TCE
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLK ;
input CLKDIV ;
input D1 ;
input D2 ;
input D3 ;
input D4 ;
input D5 ;
input D6 ;
input D7 ;
input D8 ;
input OCE ;
input RST ;
input SHIFTIN1 ;
input SHIFTIN2 ;
input T1 ;
input T2 ;
input T3 ;
input T4 ;
input TBYTEIN ;
input TCE ;
output OFB ;
output OQ ;
output SHIFTOUT1 ;
output SHIFTOUT2 ;
output TBYTEOUT ;
output TFB ;
output TQ ;
parameter DATA_RATE_OQ = "DDR";
parameter DATA_RATE_TQ = "DDR";
parameter DATA_WIDTH = 4;
parameter [0:0] INIT_OQ = 1'b0;
parameter [0:0] INIT_TQ = 1'b0;
parameter SERDES_MODE = "MASTER";
parameter [0:0] SRVAL_OQ = 1'b0;
parameter [0:0] SRVAL_TQ = 1'b0;
parameter TBYTE_CTL = "FALSE";
parameter TBYTE_SRC = "FALSE";
parameter TRISTATE_WIDTH = 4;
endmodule
//#### END MODULE DEFINITION FOR: OSERDESE2 ####

//#### BEGIN MODULE DEFINITION FOR :OUT_FIFO ###
module OUT_FIFO (
  ALMOSTEMPTY,
  ALMOSTFULL,
  EMPTY,
  FULL,
  Q0,
  Q1,
  Q2,
  Q3,
  Q4,
  Q5,
  Q6,
  Q7,
  Q8,
  Q9,

  D0,
  D1,
  D2,
  D3,
  D4,
  D5,
  D6,
  D7,
  D8,
  D9,
  RDCLK,
  RDEN,
  RESET,
  WRCLK,
  WREN
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input RDCLK ;
input RDEN ;
input RESET ;
input WRCLK ;
input WREN ;
input [7:0] D0 ;
input [7:0] D1 ;
input [7:0] D2 ;
input [7:0] D3 ;
input [7:0] D4 ;
input [7:0] D5 ;
input [7:0] D6 ;
input [7:0] D7 ;
input [7:0] D8 ;
input [7:0] D9 ;
output ALMOSTEMPTY ;
output ALMOSTFULL ;
output EMPTY ;
output FULL ;
output [3:0] Q0 ;
output [3:0] Q1 ;
output [3:0] Q2 ;
output [3:0] Q3 ;
output [3:0] Q4 ;
output [3:0] Q7 ;
output [3:0] Q8 ;
output [3:0] Q9 ;
output [7:0] Q5 ;
output [7:0] Q6 ;
parameter ALMOST_EMPTY_VALUE = 1;
parameter ALMOST_FULL_VALUE = 1;
parameter ARRAY_MODE = "ARRAY_MODE_8_X_4";
parameter OUTPUT_DISABLE = "FALSE";
parameter SYNCHRONOUS_MODE = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: OUT_FIFO ####

//#### BEGIN MODULE DEFINITION FOR :PCIE_2_0 ###
module PCIE_2_0 (
  CFGAERECRCCHECKEN,
  CFGAERECRCGENEN,
  CFGCOMMANDBUSMASTERENABLE,
  CFGCOMMANDINTERRUPTDISABLE,
  CFGCOMMANDIOENABLE,
  CFGCOMMANDMEMENABLE,
  CFGCOMMANDSERREN,
  CFGDEVCONTROL2CPLTIMEOUTDIS,
  CFGDEVCONTROL2CPLTIMEOUTVAL,
  CFGDEVCONTROLAUXPOWEREN,
  CFGDEVCONTROLCORRERRREPORTINGEN,
  CFGDEVCONTROLENABLERO,
  CFGDEVCONTROLEXTTAGEN,
  CFGDEVCONTROLFATALERRREPORTINGEN,
  CFGDEVCONTROLMAXPAYLOAD,
  CFGDEVCONTROLMAXREADREQ,
  CFGDEVCONTROLNONFATALREPORTINGEN,
  CFGDEVCONTROLNOSNOOPEN,
  CFGDEVCONTROLPHANTOMEN,
  CFGDEVCONTROLURERRREPORTINGEN,
  CFGDEVSTATUSCORRERRDETECTED,
  CFGDEVSTATUSFATALERRDETECTED,
  CFGDEVSTATUSNONFATALERRDETECTED,
  CFGDEVSTATUSURDETECTED,
  CFGDO,
  CFGERRAERHEADERLOGSETN,
  CFGERRCPLRDYN,
  CFGINTERRUPTDO,
  CFGINTERRUPTMMENABLE,
  CFGINTERRUPTMSIENABLE,
  CFGINTERRUPTMSIXENABLE,
  CFGINTERRUPTMSIXFM,
  CFGINTERRUPTRDYN,
  CFGLINKCONTROLASPMCONTROL,
  CFGLINKCONTROLAUTOBANDWIDTHINTEN,
  CFGLINKCONTROLBANDWIDTHINTEN,
  CFGLINKCONTROLCLOCKPMEN,
  CFGLINKCONTROLCOMMONCLOCK,
  CFGLINKCONTROLEXTENDEDSYNC,
  CFGLINKCONTROLHWAUTOWIDTHDIS,
  CFGLINKCONTROLLINKDISABLE,
  CFGLINKCONTROLRCB,
  CFGLINKCONTROLRETRAINLINK,
  CFGLINKSTATUSAUTOBANDWIDTHSTATUS,
  CFGLINKSTATUSBANDWITHSTATUS,
  CFGLINKSTATUSCURRENTSPEED,
  CFGLINKSTATUSDLLACTIVE,
  CFGLINKSTATUSLINKTRAINING,
  CFGLINKSTATUSNEGOTIATEDWIDTH,
  CFGMSGDATA,
  CFGMSGRECEIVED,
  CFGMSGRECEIVEDASSERTINTA,
  CFGMSGRECEIVEDASSERTINTB,
  CFGMSGRECEIVEDASSERTINTC,
  CFGMSGRECEIVEDASSERTINTD,
  CFGMSGRECEIVEDDEASSERTINTA,
  CFGMSGRECEIVEDDEASSERTINTB,
  CFGMSGRECEIVEDDEASSERTINTC,
  CFGMSGRECEIVEDDEASSERTINTD,
  CFGMSGRECEIVEDERRCOR,
  CFGMSGRECEIVEDERRFATAL,
  CFGMSGRECEIVEDERRNONFATAL,
  CFGMSGRECEIVEDPMASNAK,
  CFGMSGRECEIVEDPMETO,
  CFGMSGRECEIVEDPMETOACK,
  CFGMSGRECEIVEDPMPME,
  CFGMSGRECEIVEDSETSLOTPOWERLIMIT,
  CFGMSGRECEIVEDUNLOCK,
  CFGPCIELINKSTATE,
  CFGPMCSRPMEEN,
  CFGPMCSRPMESTATUS,
  CFGPMCSRPOWERSTATE,	 
  CFGPMRCVASREQL1N,
  CFGPMRCVENTERL1N,
  CFGPMRCVENTERL23N,
  CFGPMRCVREQACKN,
  CFGRDWRDONEN,
  CFGSLOTCONTROLELECTROMECHILCTLPULSE,
  CFGTRANSACTION,
  CFGTRANSACTIONADDR,
  CFGTRANSACTIONTYPE,
  CFGVCTCVCMAP,
  DBGSCLRA,
  DBGSCLRB,
  DBGSCLRC,
  DBGSCLRD,
  DBGSCLRE,
  DBGSCLRF,
  DBGSCLRG,
  DBGSCLRH,
  DBGSCLRI,
  DBGSCLRJ,
  DBGSCLRK,
  DBGVECA,
  DBGVECB,
  DBGVECC,
  DRPDO,
  DRPDRDY,
  LL2BADDLLPERRN,
  LL2BADTLPERRN,
  LL2PROTOCOLERRN,
  LL2REPLAYROERRN,
  LL2REPLAYTOERRN,
  LL2SUSPENDOKN,
  LL2TFCINIT1SEQN,
  LL2TFCINIT2SEQN,
  LNKCLKEN,		 
  MIMRXRADDR,
  MIMRXRCE,
  MIMRXREN,
  MIMRXWADDR,
  MIMRXWDATA,
  MIMRXWEN,
  MIMTXRADDR,
  MIMTXRCE,
  MIMTXREN,
  MIMTXWADDR,
  MIMTXWDATA,
  MIMTXWEN,
  PIPERX0POLARITY,
  PIPERX1POLARITY,
  PIPERX2POLARITY,
  PIPERX3POLARITY,
  PIPERX4POLARITY,
  PIPERX5POLARITY,
  PIPERX6POLARITY,
  PIPERX7POLARITY,
  PIPETX0CHARISK,
  PIPETX0COMPLIANCE,
  PIPETX0DATA,
  PIPETX0ELECIDLE,
  PIPETX0POWERDOWN,
  PIPETX1CHARISK,
  PIPETX1COMPLIANCE,
  PIPETX1DATA,
  PIPETX1ELECIDLE,
  PIPETX1POWERDOWN,
  PIPETX2CHARISK,
  PIPETX2COMPLIANCE,
  PIPETX2DATA,
  PIPETX2ELECIDLE,
  PIPETX2POWERDOWN,
  PIPETX3CHARISK,
  PIPETX3COMPLIANCE,
  PIPETX3DATA,
  PIPETX3ELECIDLE,
  PIPETX3POWERDOWN,
  PIPETX4CHARISK,
  PIPETX4COMPLIANCE,
  PIPETX4DATA,
  PIPETX4ELECIDLE,
  PIPETX4POWERDOWN,
  PIPETX5CHARISK,
  PIPETX5COMPLIANCE,
  PIPETX5DATA,
  PIPETX5ELECIDLE,
  PIPETX5POWERDOWN,
  PIPETX6CHARISK,
  PIPETX6COMPLIANCE,
  PIPETX6DATA,
  PIPETX6ELECIDLE,
  PIPETX6POWERDOWN,
  PIPETX7CHARISK,
  PIPETX7COMPLIANCE,
  PIPETX7DATA,
  PIPETX7ELECIDLE,
  PIPETX7POWERDOWN,
  PIPETXDEEMPH,
  PIPETXMARGIN,
  PIPETXRATE,
  PIPETXRCVRDET,
  PIPETXRESET,
  PL2LINKUPN,
  PL2RECEIVERERRN,
  PL2RECOVERYN,
  PL2RXELECIDLE,
  PL2SUSPENDOK,
  PLDBGVEC,
  PLINITIALLINKWIDTH,
  PLLANEREVERSALMODE,
  PLLINKGEN2CAP,
  PLLINKPARTNERGEN2SUPPORTED,
  PLLINKUPCFGCAP,
  PLLTSSMSTATE,
  PLPHYLNKUPN,
  PLRECEIVEDHOTRST,
  PLRXPMSTATE,
  PLSELLNKRATE,
  PLSELLNKWIDTH,
  PLTXPMSTATE,
  RECEIVEDFUNCLVLRSTN,
  TL2ASPMSUSPENDCREDITCHECKOKN,
  TL2ASPMSUSPENDREQN,
  TL2PPMSUSPENDOKN,
  TRNFCCPLD,
  TRNFCCPLH,
  TRNFCNPD,
  TRNFCNPH,
  TRNFCPD,
  TRNFCPH,
  TRNLNKUPN,
  TRNRBARHITN,
  TRNRD,
  TRNRDLLPDATA,
  TRNRDLLPSRCRDYN,
  TRNRECRCERRN,
  TRNREOFN,
  TRNRERRFWDN,
  TRNRREMN,
  TRNRSOFN,
  TRNRSRCDSCN,
  TRNRSRCRDYN,
  TRNTBUFAV,
  TRNTCFGREQN,
  TRNTDLLPDSTRDYN,
  TRNTDSTRDYN,
  TRNTERRDROPN,
  USERRSTN,
  CFGBYTEENN,
  CFGDI,
  CFGDSBUSNUMBER,
  CFGDSDEVICENUMBER,
  CFGDSFUNCTIONNUMBER,
  CFGDSN,
  CFGDWADDR,
  CFGERRACSN,
  CFGERRAERHEADERLOG,
  CFGERRCORN,
  CFGERRCPLABORTN,
  CFGERRCPLTIMEOUTN,
  CFGERRCPLUNEXPECTN,
  CFGERRECRCN,
  CFGERRLOCKEDN,
  CFGERRPOSTEDN,
  CFGERRTLPCPLHEADER,
  CFGERRURN,
  CFGINTERRUPTASSERTN,
  CFGINTERRUPTDI,
  CFGINTERRUPTN,
  CFGPMDIRECTASPML1N,
  CFGPMSENDPMACKN,
  CFGPMSENDPMETON,
  CFGPMSENDPMNAKN,
  CFGPMTURNOFFOKN,
  CFGPMWAKEN,
  CFGPORTNUMBER,
  CFGRDENN,
  CFGTRNPENDINGN,
  CFGWRENN,
  CFGWRREADONLYN,
  CFGWRRW1CASRWN,
  CMRSTN,
  CMSTICKYRSTN,
  DBGMODE,
  DBGSUBMODE,
  DLRSTN,
  DRPCLK,
  DRPDADDR,
  DRPDEN,
  DRPDI,
  DRPDWE,
  FUNCLVLRSTN,
  LL2SENDASREQL1N,
  LL2SENDENTERL1N,
  LL2SENDENTERL23N,
  LL2SUSPENDNOWN,
  LL2TLPRCVN,
  MIMRXRDATA,
  MIMTXRDATA,
  PIPECLK,
  PIPERX0CHANISALIGNED,
  PIPERX0CHARISK,
  PIPERX0DATA,
  PIPERX0ELECIDLE,
  PIPERX0PHYSTATUS,
  PIPERX0STATUS,
  PIPERX0VALID,
  PIPERX1CHANISALIGNED,
  PIPERX1CHARISK,
  PIPERX1DATA,
  PIPERX1ELECIDLE,
  PIPERX1PHYSTATUS,
  PIPERX1STATUS,
  PIPERX1VALID,
  PIPERX2CHANISALIGNED,
  PIPERX2CHARISK,
  PIPERX2DATA,
  PIPERX2ELECIDLE,
  PIPERX2PHYSTATUS,
  PIPERX2STATUS,
  PIPERX2VALID,
  PIPERX3CHANISALIGNED,
  PIPERX3CHARISK,
  PIPERX3DATA,
  PIPERX3ELECIDLE,
  PIPERX3PHYSTATUS,
  PIPERX3STATUS,
  PIPERX3VALID,
  PIPERX4CHANISALIGNED,
  PIPERX4CHARISK,
  PIPERX4DATA,
  PIPERX4ELECIDLE,
  PIPERX4PHYSTATUS,
  PIPERX4STATUS,
  PIPERX4VALID,
  PIPERX5CHANISALIGNED,
  PIPERX5CHARISK,
  PIPERX5DATA,
  PIPERX5ELECIDLE,
  PIPERX5PHYSTATUS,
  PIPERX5STATUS,
  PIPERX5VALID,
  PIPERX6CHANISALIGNED,
  PIPERX6CHARISK,
  PIPERX6DATA,
  PIPERX6ELECIDLE,
  PIPERX6PHYSTATUS,
  PIPERX6STATUS,
  PIPERX6VALID,
  PIPERX7CHANISALIGNED,
  PIPERX7CHARISK,
  PIPERX7DATA,
  PIPERX7ELECIDLE,
  PIPERX7PHYSTATUS,
  PIPERX7STATUS,
  PIPERX7VALID,
  PL2DIRECTEDLSTATE,
  PLDBGMODE,
  PLDIRECTEDLINKAUTON,
  PLDIRECTEDLINKCHANGE,
  PLDIRECTEDLINKSPEED,
  PLDIRECTEDLINKWIDTH,
  PLDOWNSTREAMDEEMPHSOURCE,
  PLRSTN,
  PLTRANSMITHOTRST,
  PLUPSTREAMPREFERDEEMPH,
  SYSRSTN,
  TL2ASPMSUSPENDCREDITCHECKN,
  TL2PPMSUSPENDREQN,
  TLRSTN,
  TRNFCSEL,
  TRNRDSTRDYN,
  TRNRNPOKN,
  TRNTCFGGNTN,
  TRNTD,
  TRNTDLLPDATA,
  TRNTDLLPSRCRDYN,
  TRNTECRCGENN,
  TRNTEOFN,
  TRNTERRFWDN,
  TRNTREMN,
  TRNTSOFN,
  TRNTSRCDSCN,
  TRNTSRCRDYN,
  TRNTSTRN,
  USERCLK
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CFGERRACSN ;
input CFGERRCORN ;
input CFGERRCPLABORTN ;
input CFGERRCPLTIMEOUTN ;
input CFGERRCPLUNEXPECTN ;
input CFGERRECRCN ;
input CFGERRLOCKEDN ;
input CFGERRPOSTEDN ;
input CFGERRURN ;
input CFGINTERRUPTASSERTN ;
input CFGINTERRUPTN ;
input CFGPMDIRECTASPML1N ;
input CFGPMSENDPMACKN ;
input CFGPMSENDPMETON ;
input CFGPMSENDPMNAKN ;
input CFGPMTURNOFFOKN ;
input CFGPMWAKEN ;
input CFGRDENN ;
input CFGTRNPENDINGN ;
input CFGWRENN ;
input CFGWRREADONLYN ;
input CFGWRRW1CASRWN ;
input CMRSTN ;
input CMSTICKYRSTN ;
input DBGSUBMODE ;
input DLRSTN ;
input DRPCLK ;
input DRPDEN ;
input DRPDWE ;
input FUNCLVLRSTN ;
input LL2SENDASREQL1N ;
input LL2SENDENTERL1N ;
input LL2SENDENTERL23N ;
input LL2SUSPENDNOWN ;
input LL2TLPRCVN ;
input PIPECLK ;
input PIPERX0CHANISALIGNED ;
input PIPERX0ELECIDLE ;
input PIPERX0PHYSTATUS ;
input PIPERX0VALID ;
input PIPERX1CHANISALIGNED ;
input PIPERX1ELECIDLE ;
input PIPERX1PHYSTATUS ;
input PIPERX1VALID ;
input PIPERX2CHANISALIGNED ;
input PIPERX2ELECIDLE ;
input PIPERX2PHYSTATUS ;
input PIPERX2VALID ;
input PIPERX3CHANISALIGNED ;
input PIPERX3ELECIDLE ;
input PIPERX3PHYSTATUS ;
input PIPERX3VALID ;
input PIPERX4CHANISALIGNED ;
input PIPERX4ELECIDLE ;
input PIPERX4PHYSTATUS ;
input PIPERX4VALID ;
input PIPERX5CHANISALIGNED ;
input PIPERX5ELECIDLE ;
input PIPERX5PHYSTATUS ;
input PIPERX5VALID ;
input PIPERX6CHANISALIGNED ;
input PIPERX6ELECIDLE ;
input PIPERX6PHYSTATUS ;
input PIPERX6VALID ;
input PIPERX7CHANISALIGNED ;
input PIPERX7ELECIDLE ;
input PIPERX7PHYSTATUS ;
input PIPERX7VALID ;
input PLDIRECTEDLINKAUTON ;
input PLDIRECTEDLINKSPEED ;
input PLDOWNSTREAMDEEMPHSOURCE ;
input PLRSTN ;
input PLTRANSMITHOTRST ;
input PLUPSTREAMPREFERDEEMPH ;
input SYSRSTN ;
input TL2ASPMSUSPENDCREDITCHECKN ;
input TL2PPMSUSPENDREQN ;
input TLRSTN ;
input TRNRDSTRDYN ;
input TRNRNPOKN ;
input TRNTCFGGNTN ;
input TRNTDLLPSRCRDYN ;
input TRNTECRCGENN ;
input TRNTEOFN ;
input TRNTERRFWDN ;
input TRNTREMN ;
input TRNTSOFN ;
input TRNTSRCDSCN ;
input TRNTSRCRDYN ;
input TRNTSTRN ;
input USERCLK ;
input [127:0] CFGERRAERHEADERLOG ;
input [15:0] DRPDI ;
input [15:0] PIPERX0DATA ;
input [15:0] PIPERX1DATA ;
input [15:0] PIPERX2DATA ;
input [15:0] PIPERX3DATA ;
input [15:0] PIPERX4DATA ;
input [15:0] PIPERX5DATA ;
input [15:0] PIPERX6DATA ;
input [15:0] PIPERX7DATA ;
input [1:0] DBGMODE ;
input [1:0] PIPERX0CHARISK ;
input [1:0] PIPERX1CHARISK ;
input [1:0] PIPERX2CHARISK ;
input [1:0] PIPERX3CHARISK ;
input [1:0] PIPERX4CHARISK ;
input [1:0] PIPERX5CHARISK ;
input [1:0] PIPERX6CHARISK ;
input [1:0] PIPERX7CHARISK ;
input [1:0] PLDIRECTEDLINKCHANGE ;
input [1:0] PLDIRECTEDLINKWIDTH ;
input [2:0] CFGDSFUNCTIONNUMBER ;
input [2:0] PIPERX0STATUS ;
input [2:0] PIPERX1STATUS ;
input [2:0] PIPERX2STATUS ;
input [2:0] PIPERX3STATUS ;
input [2:0] PIPERX4STATUS ;
input [2:0] PIPERX5STATUS ;
input [2:0] PIPERX6STATUS ;
input [2:0] PIPERX7STATUS ;
input [2:0] PLDBGMODE ;
input [2:0] TRNFCSEL ;
input [31:0] CFGDI ;
input [31:0] TRNTDLLPDATA ;
input [3:0] CFGBYTEENN ;
input [47:0] CFGERRTLPCPLHEADER ;
input [4:0] CFGDSDEVICENUMBER ;
input [4:0] PL2DIRECTEDLSTATE ;
input [63:0] CFGDSN ;
input [63:0] TRNTD ;
input [67:0] MIMRXRDATA ;
input [68:0] MIMTXRDATA ;
input [7:0] CFGDSBUSNUMBER ;
input [7:0] CFGINTERRUPTDI ;
input [7:0] CFGPORTNUMBER ;
input [8:0] DRPDADDR ;
input [9:0] CFGDWADDR ;
output CFGAERECRCCHECKEN ;
output CFGAERECRCGENEN ;
output CFGCOMMANDBUSMASTERENABLE ;
output CFGCOMMANDINTERRUPTDISABLE ;
output CFGCOMMANDIOENABLE ;
output CFGCOMMANDMEMENABLE ;
output CFGCOMMANDSERREN ;
output CFGDEVCONTROL2CPLTIMEOUTDIS ;
output CFGDEVCONTROLAUXPOWEREN ;
output CFGDEVCONTROLCORRERRREPORTINGEN ;
output CFGDEVCONTROLENABLERO ;
output CFGDEVCONTROLEXTTAGEN ;
output CFGDEVCONTROLFATALERRREPORTINGEN ;
output CFGDEVCONTROLNONFATALREPORTINGEN ;
output CFGDEVCONTROLNOSNOOPEN ;
output CFGDEVCONTROLPHANTOMEN ;
output CFGDEVCONTROLURERRREPORTINGEN ;
output CFGDEVSTATUSCORRERRDETECTED ;
output CFGDEVSTATUSFATALERRDETECTED ;
output CFGDEVSTATUSNONFATALERRDETECTED ;
output CFGDEVSTATUSURDETECTED ;
output CFGERRAERHEADERLOGSETN ;
output CFGERRCPLRDYN ;
output CFGINTERRUPTMSIENABLE ;
output CFGINTERRUPTMSIXENABLE ;
output CFGINTERRUPTMSIXFM ;
output CFGINTERRUPTRDYN ;
output CFGLINKCONTROLAUTOBANDWIDTHINTEN ;
output CFGLINKCONTROLBANDWIDTHINTEN ;
output CFGLINKCONTROLCLOCKPMEN ;
output CFGLINKCONTROLCOMMONCLOCK ;
output CFGLINKCONTROLEXTENDEDSYNC ;
output CFGLINKCONTROLHWAUTOWIDTHDIS ;
output CFGLINKCONTROLLINKDISABLE ;
output CFGLINKCONTROLRCB ;
output CFGLINKCONTROLRETRAINLINK ;
output CFGLINKSTATUSAUTOBANDWIDTHSTATUS ;
output CFGLINKSTATUSBANDWITHSTATUS ;
output CFGLINKSTATUSDLLACTIVE ;
output CFGLINKSTATUSLINKTRAINING ;
output CFGMSGRECEIVED ;
output CFGMSGRECEIVEDASSERTINTA ;
output CFGMSGRECEIVEDASSERTINTB ;
output CFGMSGRECEIVEDASSERTINTC ;
output CFGMSGRECEIVEDASSERTINTD ;
output CFGMSGRECEIVEDDEASSERTINTA ;
output CFGMSGRECEIVEDDEASSERTINTB ;
output CFGMSGRECEIVEDDEASSERTINTC ;
output CFGMSGRECEIVEDDEASSERTINTD ;
output CFGMSGRECEIVEDERRCOR ;
output CFGMSGRECEIVEDERRFATAL ;
output CFGMSGRECEIVEDERRNONFATAL ;
output CFGMSGRECEIVEDPMASNAK ;
output CFGMSGRECEIVEDPMETO ;
output CFGMSGRECEIVEDPMETOACK ;
output CFGMSGRECEIVEDPMPME ;
output CFGMSGRECEIVEDSETSLOTPOWERLIMIT ;
output CFGMSGRECEIVEDUNLOCK ;
output CFGPMCSRPMEEN ;
output CFGPMCSRPMESTATUS ;
output CFGPMRCVASREQL1N ;
output CFGPMRCVENTERL1N ;
output CFGPMRCVENTERL23N ;
output CFGPMRCVREQACKN ;
output CFGRDWRDONEN ;
output CFGSLOTCONTROLELECTROMECHILCTLPULSE ;
output CFGTRANSACTION ;
output CFGTRANSACTIONTYPE ;
output DBGSCLRA ;
output DBGSCLRB ;
output DBGSCLRC ;
output DBGSCLRD ;
output DBGSCLRE ;
output DBGSCLRF ;
output DBGSCLRG ;
output DBGSCLRH ;
output DBGSCLRI ;
output DBGSCLRJ ;
output DBGSCLRK ;
output DRPDRDY ;
output LL2BADDLLPERRN ;
output LL2BADTLPERRN ;
output LL2PROTOCOLERRN ;
output LL2REPLAYROERRN ;
output LL2REPLAYTOERRN ;
output LL2SUSPENDOKN ;
output LL2TFCINIT1SEQN ;
output LL2TFCINIT2SEQN ;
output LNKCLKEN ;
output MIMRXRCE ;
output MIMRXREN ;
output MIMRXWEN ;
output MIMTXRCE ;
output MIMTXREN ;
output MIMTXWEN ;
output PIPERX0POLARITY ;
output PIPERX1POLARITY ;
output PIPERX2POLARITY ;
output PIPERX3POLARITY ;
output PIPERX4POLARITY ;
output PIPERX5POLARITY ;
output PIPERX6POLARITY ;
output PIPERX7POLARITY ;
output PIPETX0COMPLIANCE ;
output PIPETX0ELECIDLE ;
output PIPETX1COMPLIANCE ;
output PIPETX1ELECIDLE ;
output PIPETX2COMPLIANCE ;
output PIPETX2ELECIDLE ;
output PIPETX3COMPLIANCE ;
output PIPETX3ELECIDLE ;
output PIPETX4COMPLIANCE ;
output PIPETX4ELECIDLE ;
output PIPETX5COMPLIANCE ;
output PIPETX5ELECIDLE ;
output PIPETX6COMPLIANCE ;
output PIPETX6ELECIDLE ;
output PIPETX7COMPLIANCE ;
output PIPETX7ELECIDLE ;
output PIPETXDEEMPH ;
output PIPETXRATE ;
output PIPETXRCVRDET ;
output PIPETXRESET ;
output PL2LINKUPN ;
output PL2RECEIVERERRN ;
output PL2RECOVERYN ;
output PL2RXELECIDLE ;
output PL2SUSPENDOK ;
output PLLINKGEN2CAP ;
output PLLINKPARTNERGEN2SUPPORTED ;
output PLLINKUPCFGCAP ;
output PLPHYLNKUPN ;
output PLRECEIVEDHOTRST ;
output PLSELLNKRATE ;
output RECEIVEDFUNCLVLRSTN ;
output TL2ASPMSUSPENDCREDITCHECKOKN ;
output TL2ASPMSUSPENDREQN ;
output TL2PPMSUSPENDOKN ;
output TRNLNKUPN ;
output TRNRDLLPSRCRDYN ;
output TRNRECRCERRN ;
output TRNREOFN ;
output TRNRERRFWDN ;
output TRNRREMN ;
output TRNRSOFN ;
output TRNRSRCDSCN ;
output TRNRSRCRDYN ;
output TRNTCFGREQN ;
output TRNTDLLPDSTRDYN ;
output TRNTDSTRDYN ;
output TRNTERRDROPN ;
output USERRSTN ;
output [11:0] DBGVECC ;
output [11:0] PLDBGVEC ;
output [11:0] TRNFCCPLD ;
output [11:0] TRNFCNPD ;
output [11:0] TRNFCPD ;
output [12:0] MIMRXRADDR ;
output [12:0] MIMRXWADDR ;
output [12:0] MIMTXRADDR ;
output [12:0] MIMTXWADDR ;
output [15:0] CFGMSGDATA ;
output [15:0] DRPDO ;
output [15:0] PIPETX0DATA ;
output [15:0] PIPETX1DATA ;
output [15:0] PIPETX2DATA ;
output [15:0] PIPETX3DATA ;
output [15:0] PIPETX4DATA ;
output [15:0] PIPETX5DATA ;
output [15:0] PIPETX6DATA ;
output [15:0] PIPETX7DATA ;
output [1:0] CFGLINKCONTROLASPMCONTROL ;
output [1:0] CFGLINKSTATUSCURRENTSPEED ;
output [1:0] CFGPMCSRPOWERSTATE ;
output [1:0] PIPETX0CHARISK ;
output [1:0] PIPETX0POWERDOWN ;
output [1:0] PIPETX1CHARISK ;
output [1:0] PIPETX1POWERDOWN ;
output [1:0] PIPETX2CHARISK ;
output [1:0] PIPETX2POWERDOWN ;
output [1:0] PIPETX3CHARISK ;
output [1:0] PIPETX3POWERDOWN ;
output [1:0] PIPETX4CHARISK ;
output [1:0] PIPETX4POWERDOWN ;
output [1:0] PIPETX5CHARISK ;
output [1:0] PIPETX5POWERDOWN ;
output [1:0] PIPETX6CHARISK ;
output [1:0] PIPETX6POWERDOWN ;
output [1:0] PIPETX7CHARISK ;
output [1:0] PIPETX7POWERDOWN ;
output [1:0] PLLANEREVERSALMODE ;
output [1:0] PLRXPMSTATE ;
output [1:0] PLSELLNKWIDTH ;
output [2:0] CFGDEVCONTROLMAXPAYLOAD ;
output [2:0] CFGDEVCONTROLMAXREADREQ ;
output [2:0] CFGINTERRUPTMMENABLE ;
output [2:0] CFGPCIELINKSTATE ;
output [2:0] PIPETXMARGIN ;
output [2:0] PLINITIALLINKWIDTH ;
output [2:0] PLTXPMSTATE ;
output [31:0] CFGDO ;
output [31:0] TRNRDLLPDATA ;
output [3:0] CFGDEVCONTROL2CPLTIMEOUTVAL ;
output [3:0] CFGLINKSTATUSNEGOTIATEDWIDTH ;
output [5:0] PLLTSSMSTATE ;
output [5:0] TRNTBUFAV ;
output [63:0] DBGVECA ;
output [63:0] DBGVECB ;
output [63:0] TRNRD ;
output [67:0] MIMRXWDATA ;
output [68:0] MIMTXWDATA ;
output [6:0] CFGTRANSACTIONADDR ;
output [6:0] CFGVCTCVCMAP ;
output [6:0] TRNRBARHITN ;
output [7:0] CFGINTERRUPTDO ;
output [7:0] TRNFCCPLH ;
output [7:0] TRNFCNPH ;
output [7:0] TRNFCPH ;
parameter [11:0] AER_BASE_PTR = 12'h128;
parameter AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
parameter AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
parameter [15:0] AER_CAP_ID = 16'h0001;
parameter [4:0] AER_CAP_INT_MSG_NUM_MSI = 5'h0A;
parameter [4:0] AER_CAP_INT_MSG_NUM_MSIX = 5'h15;
parameter [11:0] AER_CAP_NEXTPTR = 12'h160;
parameter AER_CAP_ON = "FALSE";
parameter AER_CAP_PERMIT_ROOTERR_UPDATE = "TRUE";
parameter [3:0] AER_CAP_VERSION = 4'h1;
parameter ALLOW_X8_GEN2 = "FALSE";
parameter [31:0] BAR0 = 32'hFFFFFF00;
parameter [31:0] BAR1 = 32'hFFFF0000;
parameter [31:0] BAR2 = 32'hFFFF000C;
parameter [31:0] BAR3 = 32'hFFFFFFFF;
parameter [31:0] BAR4 = 32'h00000000;
parameter [31:0] BAR5 = 32'h00000000;
parameter [7:0] CAPABILITIES_PTR = 8'h40;
parameter [31:0] CARDBUS_CIS_POINTER = 32'h00000000;
parameter [23:0] CLASS_CODE = 24'h000000;
parameter CMD_INTX_IMPLEMENTED = "TRUE";
parameter CPL_TIMEOUT_DISABLE_SUPPORTED = "FALSE";
parameter [3:0] CPL_TIMEOUT_RANGES_SUPPORTED = 4'h0;
parameter [6:0] CRM_MODULE_RSTS = 7'h00;
parameter [15:0] DEVICE_ID = 16'h0007;
parameter DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE = "TRUE";
parameter DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE = "TRUE";
parameter DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
parameter DEV_CAP_ENDPOINT_L1_LATENCY = 0;
parameter DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
parameter DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "FALSE";
parameter DEV_CAP_MAX_PAYLOAD_SUPPORTED = 2;
parameter DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT = 0;
parameter DEV_CAP_ROLE_BASED_ERROR = "TRUE";
parameter DEV_CAP_RSVD_14_12 = 0;
parameter DEV_CAP_RSVD_17_16 = 0;
parameter DEV_CAP_RSVD_31_29 = 0;
parameter DEV_CONTROL_AUX_POWER_SUPPORTED = "FALSE";
parameter DISABLE_ASPM_L1_TIMER = "FALSE";
parameter DISABLE_BAR_FILTERING = "FALSE";
parameter DISABLE_ID_CHECK = "FALSE";
parameter DISABLE_LANE_REVERSAL = "FALSE";
parameter DISABLE_RX_TC_FILTER = "FALSE";
parameter DISABLE_SCRAMBLING = "FALSE";
parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
parameter [11:0] DSN_BASE_PTR = 12'h100;
parameter [15:0] DSN_CAP_ID = 16'h0003;
parameter [11:0] DSN_CAP_NEXTPTR = 12'h000;
parameter DSN_CAP_ON = "TRUE";
parameter [3:0] DSN_CAP_VERSION = 4'h1;
parameter [10:0] ENABLE_MSG_ROUTE = 11'h000;
parameter ENABLE_RX_TD_ECRC_TRIM = "FALSE";
parameter ENTER_RVRY_EI_L0 = "TRUE";
parameter EXIT_LOOPBACK_ON_EI = "TRUE";
parameter [31:0] EXPANSION_ROM = 32'hFFFFF001;
parameter [5:0] EXT_CFG_CAP_PTR = 6'h3F;
parameter [9:0] EXT_CFG_XP_CAP_PTR = 10'h3FF;
parameter [7:0] HEADER_TYPE = 8'h00;
parameter [4:0] INFER_EI = 5'h00;
parameter [7:0] INTERRUPT_PIN = 8'h01;
parameter IS_SWITCH = "FALSE";
parameter [9:0] LAST_CONFIG_DWORD = 10'h042;
parameter LINK_CAP_ASPM_SUPPORT = 1;
parameter LINK_CAP_CLOCK_POWER_MANAGEMENT = "FALSE";
parameter LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP = "FALSE";
parameter LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
parameter LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
parameter LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
parameter LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
parameter LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
parameter LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
parameter LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
parameter LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
parameter LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP = "FALSE";
parameter [3:0] LINK_CAP_MAX_LINK_SPEED = 4'h1;
parameter [5:0] LINK_CAP_MAX_LINK_WIDTH = 6'h08;
parameter LINK_CAP_RSVD_23_22 = 0;
parameter LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE = "FALSE";
parameter LINK_CONTROL_RCB = 0;
parameter LINK_CTRL2_DEEMPHASIS = "FALSE";
parameter LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE = "FALSE";
parameter [3:0] LINK_CTRL2_TARGET_LINK_SPEED = 4'h2;
parameter LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
parameter [14:0] LL_ACK_TIMEOUT = 15'h0000;
parameter LL_ACK_TIMEOUT_EN = "FALSE";
parameter LL_ACK_TIMEOUT_FUNC = 0;
parameter [14:0] LL_REPLAY_TIMEOUT = 15'h0000;
parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
parameter LL_REPLAY_TIMEOUT_FUNC = 0;
parameter [5:0] LTSSM_MAX_LINK_WIDTH = 6'h01;
parameter [7:0] MSIX_BASE_PTR = 8'h9C;
parameter [7:0] MSIX_CAP_ID = 8'h11;
parameter [7:0] MSIX_CAP_NEXTPTR = 8'h00;
parameter MSIX_CAP_ON = "FALSE";
parameter MSIX_CAP_PBA_BIR = 0;
parameter [28:0] MSIX_CAP_PBA_OFFSET = 29'h00000050;
parameter MSIX_CAP_TABLE_BIR = 0;
parameter [28:0] MSIX_CAP_TABLE_OFFSET = 29'h00000040;
parameter [10:0] MSIX_CAP_TABLE_SIZE = 11'h000;
parameter [7:0] MSI_BASE_PTR = 8'h48;
parameter MSI_CAP_64_BIT_ADDR_CAPABLE = "TRUE";
parameter [7:0] MSI_CAP_ID = 8'h05;
parameter MSI_CAP_MULTIMSGCAP = 0;
parameter MSI_CAP_MULTIMSG_EXTENSION = 0;
parameter [7:0] MSI_CAP_NEXTPTR = 8'h60;
parameter MSI_CAP_ON = "FALSE";
parameter MSI_CAP_PER_VECTOR_MASKING_CAPABLE = "TRUE";
parameter N_FTS_COMCLK_GEN1 = 255;
parameter N_FTS_COMCLK_GEN2 = 255;
parameter N_FTS_GEN1 = 255;
parameter N_FTS_GEN2 = 255;
parameter [7:0] PCIE_BASE_PTR = 8'h60;
parameter [7:0] PCIE_CAP_CAPABILITY_ID = 8'h10;
parameter [3:0] PCIE_CAP_CAPABILITY_VERSION = 4'h2;
parameter [3:0] PCIE_CAP_DEVICE_PORT_TYPE = 4'h0;
parameter [4:0] PCIE_CAP_INT_MSG_NUM = 5'h00;
parameter [7:0] PCIE_CAP_NEXTPTR = 8'h00;
parameter PCIE_CAP_ON = "TRUE";
parameter PCIE_CAP_RSVD_15_14 = 0;
parameter PCIE_CAP_SLOT_IMPLEMENTED = "FALSE";
parameter PCIE_REVISION = 2;
parameter PGL0_LANE = 0;
parameter PGL1_LANE = 1;
parameter PGL2_LANE = 2;
parameter PGL3_LANE = 3;
parameter PGL4_LANE = 4;
parameter PGL5_LANE = 5;
parameter PGL6_LANE = 6;
parameter PGL7_LANE = 7;
parameter PL_AUTO_CONFIG = 0;
parameter PL_FAST_TRAIN = "FALSE";
parameter [7:0] PM_BASE_PTR = 8'h40;
parameter PM_CAP_AUXCURRENT = 0;
parameter PM_CAP_D1SUPPORT = "TRUE";
parameter PM_CAP_D2SUPPORT = "TRUE";
parameter PM_CAP_DSI = "FALSE";
parameter [7:0] PM_CAP_ID = 8'h01;
parameter [7:0] PM_CAP_NEXTPTR = 8'h48;
parameter PM_CAP_ON = "TRUE";
parameter [4:0] PM_CAP_PMESUPPORT = 5'h0F;
parameter PM_CAP_PME_CLOCK = "FALSE";
parameter PM_CAP_RSVD_04 = 0;
parameter PM_CAP_VERSION = 3;
parameter PM_CSR_B2B3 = "FALSE";
parameter PM_CSR_BPCCEN = "FALSE";
parameter PM_CSR_NOSOFTRST = "TRUE";
parameter [7:0] PM_DATA0 = 8'h01;
parameter [7:0] PM_DATA1 = 8'h01;
parameter [7:0] PM_DATA2 = 8'h01;
parameter [7:0] PM_DATA3 = 8'h01;
parameter [7:0] PM_DATA4 = 8'h01;
parameter [7:0] PM_DATA5 = 8'h01;
parameter [7:0] PM_DATA6 = 8'h01;
parameter [7:0] PM_DATA7 = 8'h01;
parameter [1:0] PM_DATA_SCALE0 = 2'h1;
parameter [1:0] PM_DATA_SCALE1 = 2'h1;
parameter [1:0] PM_DATA_SCALE2 = 2'h1;
parameter [1:0] PM_DATA_SCALE3 = 2'h1;
parameter [1:0] PM_DATA_SCALE4 = 2'h1;
parameter [1:0] PM_DATA_SCALE5 = 2'h1;
parameter [1:0] PM_DATA_SCALE6 = 2'h1;
parameter [1:0] PM_DATA_SCALE7 = 2'h1;
parameter RECRC_CHK = 0;
parameter RECRC_CHK_TRIM = "FALSE";
parameter [7:0] REVISION_ID = 8'h00;
parameter ROOT_CAP_CRS_SW_VISIBILITY = "FALSE";
parameter SELECT_DLL_IF = "FALSE";
parameter SIM_VERSION = "1.0";
parameter SLOT_CAP_ATT_BUTTON_PRESENT = "FALSE";
parameter SLOT_CAP_ATT_INDICATOR_PRESENT = "FALSE";
parameter SLOT_CAP_ELEC_INTERLOCK_PRESENT = "FALSE";
parameter SLOT_CAP_HOTPLUG_CAPABLE = "FALSE";
parameter SLOT_CAP_HOTPLUG_SURPRISE = "FALSE";
parameter SLOT_CAP_MRL_SENSOR_PRESENT = "FALSE";
parameter SLOT_CAP_NO_CMD_COMPLETED_SUPPORT = "FALSE";
parameter [12:0] SLOT_CAP_PHYSICAL_SLOT_NUM = 13'h0000;
parameter SLOT_CAP_POWER_CONTROLLER_PRESENT = "FALSE";
parameter SLOT_CAP_POWER_INDICATOR_PRESENT = "FALSE";
parameter SLOT_CAP_SLOT_POWER_LIMIT_SCALE = 0;
parameter [7:0] SLOT_CAP_SLOT_POWER_LIMIT_VALUE = 8'h00;
parameter SPARE_BIT0 = 0;
parameter SPARE_BIT1 = 0;
parameter SPARE_BIT2 = 0;
parameter SPARE_BIT3 = 0;
parameter SPARE_BIT4 = 0;
parameter SPARE_BIT5 = 0;
parameter SPARE_BIT6 = 0;
parameter SPARE_BIT7 = 0;
parameter SPARE_BIT8 = 0;
parameter [7:0] SPARE_BYTE0 = 8'h00;
parameter [7:0] SPARE_BYTE1 = 8'h00;
parameter [7:0] SPARE_BYTE2 = 8'h00;
parameter [7:0] SPARE_BYTE3 = 8'h00;
parameter [31:0] SPARE_WORD0 = 32'h00000000;
parameter [31:0] SPARE_WORD1 = 32'h00000000;
parameter [31:0] SPARE_WORD2 = 32'h00000000;
parameter [31:0] SPARE_WORD3 = 32'h00000000;
parameter [15:0] SUBSYSTEM_ID = 16'h0007;
parameter [15:0] SUBSYSTEM_VENDOR_ID = 16'h10EE;
parameter TL_RBYPASS = "FALSE";
parameter TL_RX_RAM_RADDR_LATENCY = 0;
parameter TL_RX_RAM_RDATA_LATENCY = 2;
parameter TL_RX_RAM_WRITE_LATENCY = 0;
parameter TL_TFC_DISABLE = "FALSE";
parameter TL_TX_CHECKS_DISABLE = "FALSE";
parameter TL_TX_RAM_RADDR_LATENCY = 0;
parameter TL_TX_RAM_RDATA_LATENCY = 2;
parameter TL_TX_RAM_WRITE_LATENCY = 0;
parameter UPCONFIG_CAPABLE = "TRUE";
parameter UPSTREAM_FACING = "TRUE";
parameter UR_INV_REQ = "TRUE";
parameter USER_CLK_FREQ = 3;
parameter VC0_CPL_INFINITE = "TRUE";
parameter [12:0] VC0_RX_RAM_LIMIT = 13'h03FF;
parameter VC0_TOTAL_CREDITS_CD = 127;
parameter VC0_TOTAL_CREDITS_CH = 31;
parameter VC0_TOTAL_CREDITS_NPH = 12;
parameter VC0_TOTAL_CREDITS_PD = 288;
parameter VC0_TOTAL_CREDITS_PH = 32;
parameter VC0_TX_LASTPACKET = 31;
parameter [11:0] VC_BASE_PTR = 12'h10C;
parameter [15:0] VC_CAP_ID = 16'h0002;
parameter [11:0] VC_CAP_NEXTPTR = 12'h000;
parameter VC_CAP_ON = "FALSE";
parameter VC_CAP_REJECT_SNOOP_TRANSACTIONS = "FALSE";
parameter [3:0] VC_CAP_VERSION = 4'h1;
parameter [15:0] VENDOR_ID = 16'h10EE;
parameter [11:0] VSEC_BASE_PTR = 12'h160;
parameter [15:0] VSEC_CAP_HDR_ID = 16'h1234;
parameter [11:0] VSEC_CAP_HDR_LENGTH = 12'h018;
parameter [3:0] VSEC_CAP_HDR_REVISION = 4'h1;
parameter [15:0] VSEC_CAP_ID = 16'h000B;
parameter VSEC_CAP_IS_LINK_VISIBLE = "TRUE";
parameter [11:0] VSEC_CAP_NEXTPTR = 12'h000;
parameter VSEC_CAP_ON = "FALSE";
parameter [3:0] VSEC_CAP_VERSION = 4'h1;
endmodule
//#### END MODULE DEFINITION FOR: PCIE_2_0 ####

//#### BEGIN MODULE DEFINITION FOR :PCIE_2_1 ###
module PCIE_2_1 (
  CFGAERECRCCHECKEN,
  CFGAERECRCGENEN,
  CFGAERROOTERRCORRERRRECEIVED,
  CFGAERROOTERRCORRERRREPORTINGEN,
  CFGAERROOTERRFATALERRRECEIVED,
  CFGAERROOTERRFATALERRREPORTINGEN,
  CFGAERROOTERRNONFATALERRRECEIVED,
  CFGAERROOTERRNONFATALERRREPORTINGEN,
  CFGBRIDGESERREN,
  CFGCOMMANDBUSMASTERENABLE,
  CFGCOMMANDINTERRUPTDISABLE,
  CFGCOMMANDIOENABLE,
  CFGCOMMANDMEMENABLE,
  CFGCOMMANDSERREN,
  CFGDEVCONTROL2ARIFORWARDEN,
  CFGDEVCONTROL2ATOMICEGRESSBLOCK,
  CFGDEVCONTROL2ATOMICREQUESTEREN,
  CFGDEVCONTROL2CPLTIMEOUTDIS,
  CFGDEVCONTROL2CPLTIMEOUTVAL,
  CFGDEVCONTROL2IDOCPLEN,
  CFGDEVCONTROL2IDOREQEN,
  CFGDEVCONTROL2LTREN,
  CFGDEVCONTROL2TLPPREFIXBLOCK,
  CFGDEVCONTROLAUXPOWEREN,
  CFGDEVCONTROLCORRERRREPORTINGEN,
  CFGDEVCONTROLENABLERO,
  CFGDEVCONTROLEXTTAGEN,
  CFGDEVCONTROLFATALERRREPORTINGEN,
  CFGDEVCONTROLMAXPAYLOAD,
  CFGDEVCONTROLMAXREADREQ,
  CFGDEVCONTROLNONFATALREPORTINGEN,
  CFGDEVCONTROLNOSNOOPEN,
  CFGDEVCONTROLPHANTOMEN,
  CFGDEVCONTROLURERRREPORTINGEN,
  CFGDEVSTATUSCORRERRDETECTED,
  CFGDEVSTATUSFATALERRDETECTED,
  CFGDEVSTATUSNONFATALERRDETECTED,
  CFGDEVSTATUSURDETECTED,
  CFGERRAERHEADERLOGSETN,
  CFGERRCPLRDYN,
  CFGINTERRUPTDO,
  CFGINTERRUPTMMENABLE,
  CFGINTERRUPTMSIENABLE,
  CFGINTERRUPTMSIXENABLE,
  CFGINTERRUPTMSIXFM,
  CFGINTERRUPTRDYN,
  CFGLINKCONTROLASPMCONTROL,
  CFGLINKCONTROLAUTOBANDWIDTHINTEN,
  CFGLINKCONTROLBANDWIDTHINTEN,
  CFGLINKCONTROLCLOCKPMEN,
  CFGLINKCONTROLCOMMONCLOCK,
  CFGLINKCONTROLEXTENDEDSYNC,
  CFGLINKCONTROLHWAUTOWIDTHDIS,
  CFGLINKCONTROLLINKDISABLE,
  CFGLINKCONTROLRCB,
  CFGLINKCONTROLRETRAINLINK,
  CFGLINKSTATUSAUTOBANDWIDTHSTATUS,
  CFGLINKSTATUSBANDWIDTHSTATUS,
  CFGLINKSTATUSCURRENTSPEED,
  CFGLINKSTATUSDLLACTIVE,
  CFGLINKSTATUSLINKTRAINING,
  CFGLINKSTATUSNEGOTIATEDWIDTH,
  CFGMGMTDO,
  CFGMGMTRDWRDONEN,
  CFGMSGDATA,
  CFGMSGRECEIVED,
  CFGMSGRECEIVEDASSERTINTA,
  CFGMSGRECEIVEDASSERTINTB,
  CFGMSGRECEIVEDASSERTINTC,
  CFGMSGRECEIVEDASSERTINTD,
  CFGMSGRECEIVEDDEASSERTINTA,
  CFGMSGRECEIVEDDEASSERTINTB,
  CFGMSGRECEIVEDDEASSERTINTC,
  CFGMSGRECEIVEDDEASSERTINTD,
  CFGMSGRECEIVEDERRCOR,
  CFGMSGRECEIVEDERRFATAL,
  CFGMSGRECEIVEDERRNONFATAL,
  CFGMSGRECEIVEDPMASNAK,
  CFGMSGRECEIVEDPMETO,
  CFGMSGRECEIVEDPMETOACK,
  CFGMSGRECEIVEDPMPME,
  CFGMSGRECEIVEDSETSLOTPOWERLIMIT,
  CFGMSGRECEIVEDUNLOCK,
  CFGPCIELINKSTATE,
  CFGPMCSRPMEEN,
  CFGPMCSRPMESTATUS,
  CFGPMCSRPOWERSTATE,
  CFGPMRCVASREQL1N,
  CFGPMRCVENTERL1N,
  CFGPMRCVENTERL23N,
  CFGPMRCVREQACKN,
  CFGROOTCONTROLPMEINTEN,
  CFGROOTCONTROLSYSERRCORRERREN,
  CFGROOTCONTROLSYSERRFATALERREN,
  CFGROOTCONTROLSYSERRNONFATALERREN,
  CFGSLOTCONTROLELECTROMECHILCTLPULSE,
  CFGTRANSACTION,
  CFGTRANSACTIONADDR,
  CFGTRANSACTIONTYPE,
  CFGVCTCVCMAP,
  DBGSCLRA,
  DBGSCLRB,
  DBGSCLRC,
  DBGSCLRD,
  DBGSCLRE,
  DBGSCLRF,
  DBGSCLRG,
  DBGSCLRH,
  DBGSCLRI,
  DBGSCLRJ,
  DBGSCLRK,
  DBGVECA,
  DBGVECB,
  DBGVECC,
  DRPDO,
  DRPRDY,
  LL2BADDLLPERR,
  LL2BADTLPERR,
  LL2LINKSTATUS,
  LL2PROTOCOLERR,
  LL2RECEIVERERR,
  LL2REPLAYROERR,
  LL2REPLAYTOERR,
  LL2SUSPENDOK,
  LL2TFCINIT1SEQ,
  LL2TFCINIT2SEQ,
  LL2TXIDLE,
  LNKCLKEN,
  MIMRXRADDR,
  MIMRXREN,
  MIMRXWADDR,
  MIMRXWDATA,
  MIMRXWEN,
  MIMTXRADDR,
  MIMTXREN,
  MIMTXWADDR,
  MIMTXWDATA,
  MIMTXWEN,
  PIPERX0POLARITY,
  PIPERX1POLARITY,
  PIPERX2POLARITY,
  PIPERX3POLARITY,
  PIPERX4POLARITY,
  PIPERX5POLARITY,
  PIPERX6POLARITY,
  PIPERX7POLARITY,
  PIPETX0CHARISK,
  PIPETX0COMPLIANCE,
  PIPETX0DATA,
  PIPETX0ELECIDLE,
  PIPETX0POWERDOWN,
  PIPETX1CHARISK,
  PIPETX1COMPLIANCE,
  PIPETX1DATA,
  PIPETX1ELECIDLE,
  PIPETX1POWERDOWN,
  PIPETX2CHARISK,
  PIPETX2COMPLIANCE,
  PIPETX2DATA,
  PIPETX2ELECIDLE,
  PIPETX2POWERDOWN,
  PIPETX3CHARISK,
  PIPETX3COMPLIANCE,
  PIPETX3DATA,
  PIPETX3ELECIDLE,
  PIPETX3POWERDOWN,
  PIPETX4CHARISK,
  PIPETX4COMPLIANCE,
  PIPETX4DATA,
  PIPETX4ELECIDLE,
  PIPETX4POWERDOWN,
  PIPETX5CHARISK,
  PIPETX5COMPLIANCE,
  PIPETX5DATA,
  PIPETX5ELECIDLE,
  PIPETX5POWERDOWN,
  PIPETX6CHARISK,
  PIPETX6COMPLIANCE,
  PIPETX6DATA,
  PIPETX6ELECIDLE,
  PIPETX6POWERDOWN,
  PIPETX7CHARISK,
  PIPETX7COMPLIANCE,
  PIPETX7DATA,
  PIPETX7ELECIDLE,
  PIPETX7POWERDOWN,
  PIPETXDEEMPH,
  PIPETXMARGIN,
  PIPETXRATE,
  PIPETXRCVRDET,
  PIPETXRESET,
  PL2L0REQ,
  PL2LINKUP,
  PL2RECEIVERERR,
  PL2RECOVERY,
  PL2RXELECIDLE,
  PL2RXPMSTATE,
  PL2SUSPENDOK,
  PLDBGVEC,
  PLDIRECTEDCHANGEDONE,
  PLINITIALLINKWIDTH,
  PLLANEREVERSALMODE,
  PLLINKGEN2CAP,
  PLLINKPARTNERGEN2SUPPORTED,
  PLLINKUPCFGCAP,
  PLLTSSMSTATE,
  PLPHYLNKUPN,
  PLRECEIVEDHOTRST,
  PLRXPMSTATE,
  PLSELLNKRATE,
  PLSELLNKWIDTH,
  PLTXPMSTATE,
  RECEIVEDFUNCLVLRSTN,
  TL2ASPMSUSPENDCREDITCHECKOK,
  TL2ASPMSUSPENDREQ,
  TL2ERRFCPE,
  TL2ERRHDR,
  TL2ERRMALFORMED,
  TL2ERRRXOVERFLOW,
  TL2PPMSUSPENDOK,
  TRNFCCPLD,
  TRNFCCPLH,
  TRNFCNPD,
  TRNFCNPH,
  TRNFCPD,
  TRNFCPH,
  TRNLNKUP,
  TRNRBARHIT,
  TRNRD,
  TRNRDLLPDATA,
  TRNRDLLPSRCRDY,
  TRNRECRCERR,
  TRNREOF,
  TRNRERRFWD,
  TRNRREM,
  TRNRSOF,
  TRNRSRCDSC,
  TRNRSRCRDY,
  TRNTBUFAV,
  TRNTCFGREQ,
  TRNTDLLPDSTRDY,
  TRNTDSTRDY,
  TRNTERRDROP,
  USERRSTN,

  CFGAERINTERRUPTMSGNUM,
  CFGDEVID,
  CFGDSBUSNUMBER,
  CFGDSDEVICENUMBER,
  CFGDSFUNCTIONNUMBER,
  CFGDSN,
  CFGERRACSN,
  CFGERRAERHEADERLOG,
  CFGERRATOMICEGRESSBLOCKEDN,
  CFGERRCORN,
  CFGERRCPLABORTN,
  CFGERRCPLTIMEOUTN,
  CFGERRCPLUNEXPECTN,
  CFGERRECRCN,
  CFGERRINTERNALCORN,
  CFGERRINTERNALUNCORN,
  CFGERRLOCKEDN,
  CFGERRMALFORMEDN,
  CFGERRMCBLOCKEDN,
  CFGERRNORECOVERYN,
  CFGERRPOISONEDN,
  CFGERRPOSTEDN,
  CFGERRTLPCPLHEADER,
  CFGERRURN,
  CFGFORCECOMMONCLOCKOFF,
  CFGFORCEEXTENDEDSYNCON,
  CFGFORCEMPS,
  CFGINTERRUPTASSERTN,
  CFGINTERRUPTDI,
  CFGINTERRUPTN,
  CFGINTERRUPTSTATN,
  CFGMGMTBYTEENN,
  CFGMGMTDI,
  CFGMGMTDWADDR,
  CFGMGMTRDENN,
  CFGMGMTWRENN,
  CFGMGMTWRREADONLYN,
  CFGMGMTWRRW1CASRWN,
  CFGPCIECAPINTERRUPTMSGNUM,
  CFGPMFORCESTATE,
  CFGPMFORCESTATEENN,
  CFGPMHALTASPML0SN,
  CFGPMHALTASPML1N,
  CFGPMSENDPMETON,
  CFGPMTURNOFFOKN,
  CFGPMWAKEN,
  CFGPORTNUMBER,
  CFGREVID,
  CFGSUBSYSID,
  CFGSUBSYSVENDID,
  CFGTRNPENDINGN,
  CFGVENDID,
  CMRSTN,
  CMSTICKYRSTN,
  DBGMODE,
  DBGSUBMODE,
  DLRSTN,
  DRPADDR,
  DRPCLK,
  DRPDI,
  DRPEN,
  DRPWE,
  FUNCLVLRSTN,
  LL2SENDASREQL1,
  LL2SENDENTERL1,
  LL2SENDENTERL23,
  LL2SENDPMACK,
  LL2SUSPENDNOW,
  LL2TLPRCV,
  MIMRXRDATA,
  MIMTXRDATA,
  PIPECLK,
  PIPERX0CHANISALIGNED,
  PIPERX0CHARISK,
  PIPERX0DATA,
  PIPERX0ELECIDLE,
  PIPERX0PHYSTATUS,
  PIPERX0STATUS,
  PIPERX0VALID,
  PIPERX1CHANISALIGNED,
  PIPERX1CHARISK,
  PIPERX1DATA,
  PIPERX1ELECIDLE,
  PIPERX1PHYSTATUS,
  PIPERX1STATUS,
  PIPERX1VALID,
  PIPERX2CHANISALIGNED,
  PIPERX2CHARISK,
  PIPERX2DATA,
  PIPERX2ELECIDLE,
  PIPERX2PHYSTATUS,
  PIPERX2STATUS,
  PIPERX2VALID,
  PIPERX3CHANISALIGNED,
  PIPERX3CHARISK,
  PIPERX3DATA,
  PIPERX3ELECIDLE,
  PIPERX3PHYSTATUS,
  PIPERX3STATUS,
  PIPERX3VALID,
  PIPERX4CHANISALIGNED,
  PIPERX4CHARISK,
  PIPERX4DATA,
  PIPERX4ELECIDLE,
  PIPERX4PHYSTATUS,
  PIPERX4STATUS,
  PIPERX4VALID,
  PIPERX5CHANISALIGNED,
  PIPERX5CHARISK,
  PIPERX5DATA,
  PIPERX5ELECIDLE,
  PIPERX5PHYSTATUS,
  PIPERX5STATUS,
  PIPERX5VALID,
  PIPERX6CHANISALIGNED,
  PIPERX6CHARISK,
  PIPERX6DATA,
  PIPERX6ELECIDLE,
  PIPERX6PHYSTATUS,
  PIPERX6STATUS,
  PIPERX6VALID,
  PIPERX7CHANISALIGNED,
  PIPERX7CHARISK,
  PIPERX7DATA,
  PIPERX7ELECIDLE,
  PIPERX7PHYSTATUS,
  PIPERX7STATUS,
  PIPERX7VALID,
  PL2DIRECTEDLSTATE,
  PLDBGMODE,
  PLDIRECTEDLINKAUTON,
  PLDIRECTEDLINKCHANGE,
  PLDIRECTEDLINKSPEED,
  PLDIRECTEDLINKWIDTH,
  PLDIRECTEDLTSSMNEW,
  PLDIRECTEDLTSSMNEWVLD,
  PLDIRECTEDLTSSMSTALL,
  PLDOWNSTREAMDEEMPHSOURCE,
  PLRSTN,
  PLTRANSMITHOTRST,
  PLUPSTREAMPREFERDEEMPH,
  SYSRSTN,
  TL2ASPMSUSPENDCREDITCHECK,
  TL2PPMSUSPENDREQ,
  TLRSTN,
  TRNFCSEL,
  TRNRDSTRDY,
  TRNRFCPRET,
  TRNRNPOK,
  TRNRNPREQ,
  TRNTCFGGNT,
  TRNTD,
  TRNTDLLPDATA,
  TRNTDLLPSRCRDY,
  TRNTECRCGEN,
  TRNTEOF,
  TRNTERRFWD,
  TRNTREM,
  TRNTSOF,
  TRNTSRCDSC,
  TRNTSRCRDY,
  TRNTSTR,
  USERCLK,
  USERCLK2
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CFGERRACSN ;
input CFGERRATOMICEGRESSBLOCKEDN ;
input CFGERRCORN ;
input CFGERRCPLABORTN ;
input CFGERRCPLTIMEOUTN ;
input CFGERRCPLUNEXPECTN ;
input CFGERRECRCN ;
input CFGERRINTERNALCORN ;
input CFGERRINTERNALUNCORN ;
input CFGERRLOCKEDN ;
input CFGERRMALFORMEDN ;
input CFGERRMCBLOCKEDN ;
input CFGERRNORECOVERYN ;
input CFGERRPOISONEDN ;
input CFGERRPOSTEDN ;
input CFGERRURN ;
input CFGFORCECOMMONCLOCKOFF ;
input CFGFORCEEXTENDEDSYNCON ;
input CFGINTERRUPTASSERTN ;
input CFGINTERRUPTN ;
input CFGINTERRUPTSTATN ;
input CFGMGMTRDENN ;
input CFGMGMTWRENN ;
input CFGMGMTWRREADONLYN ;
input CFGMGMTWRRW1CASRWN ;
input CFGPMFORCESTATEENN ;
input CFGPMHALTASPML0SN ;
input CFGPMHALTASPML1N ;
input CFGPMSENDPMETON ;
input CFGPMTURNOFFOKN ;
input CFGPMWAKEN ;
input CFGTRNPENDINGN ;
input CMRSTN ;
input CMSTICKYRSTN ;
input DBGSUBMODE ;
input DLRSTN ;
input DRPCLK ;
input DRPEN ;
input DRPWE ;
input FUNCLVLRSTN ;
input LL2SENDASREQL1 ;
input LL2SENDENTERL1 ;
input LL2SENDENTERL23 ;
input LL2SENDPMACK ;
input LL2SUSPENDNOW ;
input LL2TLPRCV ;
input PIPECLK ;
input PIPERX0CHANISALIGNED ;
input PIPERX0ELECIDLE ;
input PIPERX0PHYSTATUS ;
input PIPERX0VALID ;
input PIPERX1CHANISALIGNED ;
input PIPERX1ELECIDLE ;
input PIPERX1PHYSTATUS ;
input PIPERX1VALID ;
input PIPERX2CHANISALIGNED ;
input PIPERX2ELECIDLE ;
input PIPERX2PHYSTATUS ;
input PIPERX2VALID ;
input PIPERX3CHANISALIGNED ;
input PIPERX3ELECIDLE ;
input PIPERX3PHYSTATUS ;
input PIPERX3VALID ;
input PIPERX4CHANISALIGNED ;
input PIPERX4ELECIDLE ;
input PIPERX4PHYSTATUS ;
input PIPERX4VALID ;
input PIPERX5CHANISALIGNED ;
input PIPERX5ELECIDLE ;
input PIPERX5PHYSTATUS ;
input PIPERX5VALID ;
input PIPERX6CHANISALIGNED ;
input PIPERX6ELECIDLE ;
input PIPERX6PHYSTATUS ;
input PIPERX6VALID ;
input PIPERX7CHANISALIGNED ;
input PIPERX7ELECIDLE ;
input PIPERX7PHYSTATUS ;
input PIPERX7VALID ;
input PLDIRECTEDLINKAUTON ;
input PLDIRECTEDLINKSPEED ;
input PLDIRECTEDLTSSMNEWVLD ;
input PLDIRECTEDLTSSMSTALL ;
input PLDOWNSTREAMDEEMPHSOURCE ;
input PLRSTN ;
input PLTRANSMITHOTRST ;
input PLUPSTREAMPREFERDEEMPH ;
input SYSRSTN ;
input TL2ASPMSUSPENDCREDITCHECK ;
input TL2PPMSUSPENDREQ ;
input TLRSTN ;
input TRNRDSTRDY ;
input TRNRFCPRET ;
input TRNRNPOK ;
input TRNRNPREQ ;
input TRNTCFGGNT ;
input TRNTDLLPSRCRDY ;
input TRNTECRCGEN ;
input TRNTEOF ;
input TRNTERRFWD ;
input TRNTSOF ;
input TRNTSRCDSC ;
input TRNTSRCRDY ;
input TRNTSTR ;
input USERCLK2 ;
input USERCLK ;
input [127:0] CFGERRAERHEADERLOG ;
input [127:0] TRNTD ;
input [15:0] CFGDEVID ;
input [15:0] CFGSUBSYSID ;
input [15:0] CFGSUBSYSVENDID ;
input [15:0] CFGVENDID ;
input [15:0] DRPDI ;
input [15:0] PIPERX0DATA ;
input [15:0] PIPERX1DATA ;
input [15:0] PIPERX2DATA ;
input [15:0] PIPERX3DATA ;
input [15:0] PIPERX4DATA ;
input [15:0] PIPERX5DATA ;
input [15:0] PIPERX6DATA ;
input [15:0] PIPERX7DATA ;
input [1:0] CFGPMFORCESTATE ;
input [1:0] DBGMODE ;
input [1:0] PIPERX0CHARISK ;
input [1:0] PIPERX1CHARISK ;
input [1:0] PIPERX2CHARISK ;
input [1:0] PIPERX3CHARISK ;
input [1:0] PIPERX4CHARISK ;
input [1:0] PIPERX5CHARISK ;
input [1:0] PIPERX6CHARISK ;
input [1:0] PIPERX7CHARISK ;
input [1:0] PLDIRECTEDLINKCHANGE ;
input [1:0] PLDIRECTEDLINKWIDTH ;
input [1:0] TRNTREM ;
input [2:0] CFGDSFUNCTIONNUMBER ;
input [2:0] CFGFORCEMPS ;
input [2:0] PIPERX0STATUS ;
input [2:0] PIPERX1STATUS ;
input [2:0] PIPERX2STATUS ;
input [2:0] PIPERX3STATUS ;
input [2:0] PIPERX4STATUS ;
input [2:0] PIPERX5STATUS ;
input [2:0] PIPERX6STATUS ;
input [2:0] PIPERX7STATUS ;
input [2:0] PLDBGMODE ;
input [2:0] TRNFCSEL ;
input [31:0] CFGMGMTDI ;
input [31:0] TRNTDLLPDATA ;
input [3:0] CFGMGMTBYTEENN ;
input [47:0] CFGERRTLPCPLHEADER ;
input [4:0] CFGAERINTERRUPTMSGNUM ;
input [4:0] CFGDSDEVICENUMBER ;
input [4:0] CFGPCIECAPINTERRUPTMSGNUM ;
input [4:0] PL2DIRECTEDLSTATE ;
input [5:0] PLDIRECTEDLTSSMNEW ;
input [63:0] CFGDSN ;
input [67:0] MIMRXRDATA ;
input [68:0] MIMTXRDATA ;
input [7:0] CFGDSBUSNUMBER ;
input [7:0] CFGINTERRUPTDI ;
input [7:0] CFGPORTNUMBER ;
input [7:0] CFGREVID ;
input [8:0] DRPADDR ;
input [9:0] CFGMGMTDWADDR ;
output CFGAERECRCCHECKEN ;
output CFGAERECRCGENEN ;
output CFGAERROOTERRCORRERRRECEIVED ;
output CFGAERROOTERRCORRERRREPORTINGEN ;
output CFGAERROOTERRFATALERRRECEIVED ;
output CFGAERROOTERRFATALERRREPORTINGEN ;
output CFGAERROOTERRNONFATALERRRECEIVED ;
output CFGAERROOTERRNONFATALERRREPORTINGEN ;
output CFGBRIDGESERREN ;
output CFGCOMMANDBUSMASTERENABLE ;
output CFGCOMMANDINTERRUPTDISABLE ;
output CFGCOMMANDIOENABLE ;
output CFGCOMMANDMEMENABLE ;
output CFGCOMMANDSERREN ;
output CFGDEVCONTROL2ARIFORWARDEN ;
output CFGDEVCONTROL2ATOMICEGRESSBLOCK ;
output CFGDEVCONTROL2ATOMICREQUESTEREN ;
output CFGDEVCONTROL2CPLTIMEOUTDIS ;
output CFGDEVCONTROL2IDOCPLEN ;
output CFGDEVCONTROL2IDOREQEN ;
output CFGDEVCONTROL2LTREN ;
output CFGDEVCONTROL2TLPPREFIXBLOCK ;
output CFGDEVCONTROLAUXPOWEREN ;
output CFGDEVCONTROLCORRERRREPORTINGEN ;
output CFGDEVCONTROLENABLERO ;
output CFGDEVCONTROLEXTTAGEN ;
output CFGDEVCONTROLFATALERRREPORTINGEN ;
output CFGDEVCONTROLNONFATALREPORTINGEN ;
output CFGDEVCONTROLNOSNOOPEN ;
output CFGDEVCONTROLPHANTOMEN ;
output CFGDEVCONTROLURERRREPORTINGEN ;
output CFGDEVSTATUSCORRERRDETECTED ;
output CFGDEVSTATUSFATALERRDETECTED ;
output CFGDEVSTATUSNONFATALERRDETECTED ;
output CFGDEVSTATUSURDETECTED ;
output CFGERRAERHEADERLOGSETN ;
output CFGERRCPLRDYN ;
output CFGINTERRUPTMSIENABLE ;
output CFGINTERRUPTMSIXENABLE ;
output CFGINTERRUPTMSIXFM ;
output CFGINTERRUPTRDYN ;
output CFGLINKCONTROLAUTOBANDWIDTHINTEN ;
output CFGLINKCONTROLBANDWIDTHINTEN ;
output CFGLINKCONTROLCLOCKPMEN ;
output CFGLINKCONTROLCOMMONCLOCK ;
output CFGLINKCONTROLEXTENDEDSYNC ;
output CFGLINKCONTROLHWAUTOWIDTHDIS ;
output CFGLINKCONTROLLINKDISABLE ;
output CFGLINKCONTROLRCB ;
output CFGLINKCONTROLRETRAINLINK ;
output CFGLINKSTATUSAUTOBANDWIDTHSTATUS ;
output CFGLINKSTATUSBANDWIDTHSTATUS ;
output CFGLINKSTATUSDLLACTIVE ;
output CFGLINKSTATUSLINKTRAINING ;
output CFGMGMTRDWRDONEN ;
output CFGMSGRECEIVED ;
output CFGMSGRECEIVEDASSERTINTA ;
output CFGMSGRECEIVEDASSERTINTB ;
output CFGMSGRECEIVEDASSERTINTC ;
output CFGMSGRECEIVEDASSERTINTD ;
output CFGMSGRECEIVEDDEASSERTINTA ;
output CFGMSGRECEIVEDDEASSERTINTB ;
output CFGMSGRECEIVEDDEASSERTINTC ;
output CFGMSGRECEIVEDDEASSERTINTD ;
output CFGMSGRECEIVEDERRCOR ;
output CFGMSGRECEIVEDERRFATAL ;
output CFGMSGRECEIVEDERRNONFATAL ;
output CFGMSGRECEIVEDPMASNAK ;
output CFGMSGRECEIVEDPMETO ;
output CFGMSGRECEIVEDPMETOACK ;
output CFGMSGRECEIVEDPMPME ;
output CFGMSGRECEIVEDSETSLOTPOWERLIMIT ;
output CFGMSGRECEIVEDUNLOCK ;
output CFGPMCSRPMEEN ;
output CFGPMCSRPMESTATUS ;
output CFGPMRCVASREQL1N ;
output CFGPMRCVENTERL1N ;
output CFGPMRCVENTERL23N ;
output CFGPMRCVREQACKN ;
output CFGROOTCONTROLPMEINTEN ;
output CFGROOTCONTROLSYSERRCORRERREN ;
output CFGROOTCONTROLSYSERRFATALERREN ;
output CFGROOTCONTROLSYSERRNONFATALERREN ;
output CFGSLOTCONTROLELECTROMECHILCTLPULSE ;
output CFGTRANSACTION ;
output CFGTRANSACTIONTYPE ;
output DBGSCLRA ;
output DBGSCLRB ;
output DBGSCLRC ;
output DBGSCLRD ;
output DBGSCLRE ;
output DBGSCLRF ;
output DBGSCLRG ;
output DBGSCLRH ;
output DBGSCLRI ;
output DBGSCLRJ ;
output DBGSCLRK ;
output DRPRDY ;
output LL2BADDLLPERR ;
output LL2BADTLPERR ;
output LL2PROTOCOLERR ;
output LL2RECEIVERERR ;
output LL2REPLAYROERR ;
output LL2REPLAYTOERR ;
output LL2SUSPENDOK ;
output LL2TFCINIT1SEQ ;
output LL2TFCINIT2SEQ ;
output LL2TXIDLE ;
output LNKCLKEN ;
output MIMRXREN ;
output MIMRXWEN ;
output MIMTXREN ;
output MIMTXWEN ;
output PIPERX0POLARITY ;
output PIPERX1POLARITY ;
output PIPERX2POLARITY ;
output PIPERX3POLARITY ;
output PIPERX4POLARITY ;
output PIPERX5POLARITY ;
output PIPERX6POLARITY ;
output PIPERX7POLARITY ;
output PIPETX0COMPLIANCE ;
output PIPETX0ELECIDLE ;
output PIPETX1COMPLIANCE ;
output PIPETX1ELECIDLE ;
output PIPETX2COMPLIANCE ;
output PIPETX2ELECIDLE ;
output PIPETX3COMPLIANCE ;
output PIPETX3ELECIDLE ;
output PIPETX4COMPLIANCE ;
output PIPETX4ELECIDLE ;
output PIPETX5COMPLIANCE ;
output PIPETX5ELECIDLE ;
output PIPETX6COMPLIANCE ;
output PIPETX6ELECIDLE ;
output PIPETX7COMPLIANCE ;
output PIPETX7ELECIDLE ;
output PIPETXDEEMPH ;
output PIPETXRATE ;
output PIPETXRCVRDET ;
output PIPETXRESET ;
output PL2L0REQ ;
output PL2LINKUP ;
output PL2RECEIVERERR ;
output PL2RECOVERY ;
output PL2RXELECIDLE ;
output PL2SUSPENDOK ;
output PLDIRECTEDCHANGEDONE ;
output PLLINKGEN2CAP ;
output PLLINKPARTNERGEN2SUPPORTED ;
output PLLINKUPCFGCAP ;
output PLPHYLNKUPN ;
output PLRECEIVEDHOTRST ;
output PLSELLNKRATE ;
output RECEIVEDFUNCLVLRSTN ;
output TL2ASPMSUSPENDCREDITCHECKOK ;
output TL2ASPMSUSPENDREQ ;
output TL2ERRFCPE ;
output TL2ERRMALFORMED ;
output TL2ERRRXOVERFLOW ;
output TL2PPMSUSPENDOK ;
output TRNLNKUP ;
output TRNRECRCERR ;
output TRNREOF ;
output TRNRERRFWD ;
output TRNRSOF ;
output TRNRSRCDSC ;
output TRNRSRCRDY ;
output TRNTCFGREQ ;
output TRNTDLLPDSTRDY ;
output TRNTERRDROP ;
output USERRSTN ;
output [11:0] DBGVECC ;
output [11:0] PLDBGVEC ;
output [11:0] TRNFCCPLD ;
output [11:0] TRNFCNPD ;
output [11:0] TRNFCPD ;
output [127:0] TRNRD ;
output [12:0] MIMRXRADDR ;
output [12:0] MIMRXWADDR ;
output [12:0] MIMTXRADDR ;
output [12:0] MIMTXWADDR ;
output [15:0] CFGMSGDATA ;
output [15:0] DRPDO ;
output [15:0] PIPETX0DATA ;
output [15:0] PIPETX1DATA ;
output [15:0] PIPETX2DATA ;
output [15:0] PIPETX3DATA ;
output [15:0] PIPETX4DATA ;
output [15:0] PIPETX5DATA ;
output [15:0] PIPETX6DATA ;
output [15:0] PIPETX7DATA ;
output [1:0] CFGLINKCONTROLASPMCONTROL ;
output [1:0] CFGLINKSTATUSCURRENTSPEED ;
output [1:0] CFGPMCSRPOWERSTATE ;
output [1:0] PIPETX0CHARISK ;
output [1:0] PIPETX0POWERDOWN ;
output [1:0] PIPETX1CHARISK ;
output [1:0] PIPETX1POWERDOWN ;
output [1:0] PIPETX2CHARISK ;
output [1:0] PIPETX2POWERDOWN ;
output [1:0] PIPETX3CHARISK ;
output [1:0] PIPETX3POWERDOWN ;
output [1:0] PIPETX4CHARISK ;
output [1:0] PIPETX4POWERDOWN ;
output [1:0] PIPETX5CHARISK ;
output [1:0] PIPETX5POWERDOWN ;
output [1:0] PIPETX6CHARISK ;
output [1:0] PIPETX6POWERDOWN ;
output [1:0] PIPETX7CHARISK ;
output [1:0] PIPETX7POWERDOWN ;
output [1:0] PL2RXPMSTATE ;
output [1:0] PLLANEREVERSALMODE ;
output [1:0] PLRXPMSTATE ;
output [1:0] PLSELLNKWIDTH ;
output [1:0] TRNRDLLPSRCRDY ;
output [1:0] TRNRREM ;
output [2:0] CFGDEVCONTROLMAXPAYLOAD ;
output [2:0] CFGDEVCONTROLMAXREADREQ ;
output [2:0] CFGINTERRUPTMMENABLE ;
output [2:0] CFGPCIELINKSTATE ;
output [2:0] PIPETXMARGIN ;
output [2:0] PLINITIALLINKWIDTH ;
output [2:0] PLTXPMSTATE ;
output [31:0] CFGMGMTDO ;
output [3:0] CFGDEVCONTROL2CPLTIMEOUTVAL ;
output [3:0] CFGLINKSTATUSNEGOTIATEDWIDTH ;
output [3:0] TRNTDSTRDY ;
output [4:0] LL2LINKSTATUS ;
output [5:0] PLLTSSMSTATE ;
output [5:0] TRNTBUFAV ;
output [63:0] DBGVECA ;
output [63:0] DBGVECB ;
output [63:0] TL2ERRHDR ;
output [63:0] TRNRDLLPDATA ;
output [67:0] MIMRXWDATA ;
output [68:0] MIMTXWDATA ;
output [6:0] CFGTRANSACTIONADDR ;
output [6:0] CFGVCTCVCMAP ;
output [7:0] CFGINTERRUPTDO ;
output [7:0] TRNFCCPLH ;
output [7:0] TRNFCNPH ;
output [7:0] TRNFCPH ;
output [7:0] TRNRBARHIT ;
parameter [11:0] AER_BASE_PTR = 12'h140;
parameter AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
parameter AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
parameter [15:0] AER_CAP_ID = 16'h0001;
parameter AER_CAP_MULTIHEADER = "FALSE";
parameter [11:0] AER_CAP_NEXTPTR = 12'h178;
parameter AER_CAP_ON = "FALSE";
parameter [23:0] AER_CAP_OPTIONAL_ERR_SUPPORT = 24'h000000;
parameter AER_CAP_PERMIT_ROOTERR_UPDATE = "TRUE";
parameter [3:0] AER_CAP_VERSION = 4'h2;
parameter ALLOW_X8_GEN2 = "FALSE";
parameter [31:0] BAR0 = 32'hFFFFFF00;
parameter [31:0] BAR1 = 32'hFFFF0000;
parameter [31:0] BAR2 = 32'hFFFF000C;
parameter [31:0] BAR3 = 32'hFFFFFFFF;
parameter [31:0] BAR4 = 32'h00000000;
parameter [31:0] BAR5 = 32'h00000000;
parameter [7:0] CAPABILITIES_PTR = 8'h40;
parameter [31:0] CARDBUS_CIS_POINTER = 32'h00000000;
parameter CFG_ECRC_ERR_CPLSTAT = 0;
parameter [23:0] CLASS_CODE = 24'h000000;
parameter CMD_INTX_IMPLEMENTED = "TRUE";
parameter CPL_TIMEOUT_DISABLE_SUPPORTED = "FALSE";
parameter [3:0] CPL_TIMEOUT_RANGES_SUPPORTED = 4'h0;
parameter [6:0] CRM_MODULE_RSTS = 7'h00;
parameter DEV_CAP2_ARI_FORWARDING_SUPPORTED = "FALSE";
parameter DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED = "FALSE";
parameter DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED = "FALSE";
parameter DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED = "FALSE";
parameter DEV_CAP2_CAS128_COMPLETER_SUPPORTED = "FALSE";
parameter DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED = "FALSE";
parameter DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED = "FALSE";
parameter DEV_CAP2_LTR_MECHANISM_SUPPORTED = "FALSE";
parameter [1:0] DEV_CAP2_MAX_ENDEND_TLP_PREFIXES = 2'h0;
parameter DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING = "FALSE";
parameter [1:0] DEV_CAP2_TPH_COMPLETER_SUPPORTED = 2'h0;
parameter DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE = "TRUE";
parameter DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE = "TRUE";
parameter DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
parameter DEV_CAP_ENDPOINT_L1_LATENCY = 0;
parameter DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
parameter DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "FALSE";
parameter DEV_CAP_MAX_PAYLOAD_SUPPORTED = 2;
parameter DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT = 0;
parameter DEV_CAP_ROLE_BASED_ERROR = "TRUE";
parameter DEV_CAP_RSVD_14_12 = 0;
parameter DEV_CAP_RSVD_17_16 = 0;
parameter DEV_CAP_RSVD_31_29 = 0;
parameter DEV_CONTROL_AUX_POWER_SUPPORTED = "FALSE";
parameter DEV_CONTROL_EXT_TAG_DEFAULT = "FALSE";
parameter DISABLE_ASPM_L1_TIMER = "FALSE";
parameter DISABLE_BAR_FILTERING = "FALSE";
parameter DISABLE_ERR_MSG = "FALSE";
parameter DISABLE_ID_CHECK = "FALSE";
parameter DISABLE_LANE_REVERSAL = "FALSE";
parameter DISABLE_LOCKED_FILTER = "FALSE";
parameter DISABLE_PPM_FILTER = "FALSE";
parameter DISABLE_RX_POISONED_RESP = "FALSE";
parameter DISABLE_RX_TC_FILTER = "FALSE";
parameter DISABLE_SCRAMBLING = "FALSE";
parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
parameter [11:0] DSN_BASE_PTR = 12'h100;
parameter [15:0] DSN_CAP_ID = 16'h0003;
parameter [11:0] DSN_CAP_NEXTPTR = 12'h10C;
parameter DSN_CAP_ON = "TRUE";
parameter [3:0] DSN_CAP_VERSION = 4'h1;
parameter [10:0] ENABLE_MSG_ROUTE = 11'h000;
parameter ENABLE_RX_TD_ECRC_TRIM = "FALSE";
parameter ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED = "FALSE";
parameter ENTER_RVRY_EI_L0 = "TRUE";
parameter EXIT_LOOPBACK_ON_EI = "TRUE";
parameter [31:0] EXPANSION_ROM = 32'hFFFFF001;
parameter [5:0] EXT_CFG_CAP_PTR = 6'h3F;
parameter [9:0] EXT_CFG_XP_CAP_PTR = 10'h3FF;
parameter [7:0] HEADER_TYPE = 8'h00;
parameter [4:0] INFER_EI = 5'h00;
parameter [7:0] INTERRUPT_PIN = 8'h01;
parameter INTERRUPT_STAT_AUTO = "TRUE";
parameter IS_SWITCH = "FALSE";
parameter [9:0] LAST_CONFIG_DWORD = 10'h3FF;
parameter LINK_CAP_ASPM_OPTIONALITY = "TRUE";
parameter LINK_CAP_ASPM_SUPPORT = 1;
parameter LINK_CAP_CLOCK_POWER_MANAGEMENT = "FALSE";
parameter LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP = "FALSE";
parameter LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
parameter LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
parameter LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
parameter LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
parameter LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
parameter LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
parameter LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
parameter LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
parameter LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP = "FALSE";
parameter [3:0] LINK_CAP_MAX_LINK_SPEED = 4'h1;
parameter [5:0] LINK_CAP_MAX_LINK_WIDTH = 6'h08;
parameter LINK_CAP_RSVD_23 = 0;
parameter LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE = "FALSE";
parameter LINK_CONTROL_RCB = 0;
parameter LINK_CTRL2_DEEMPHASIS = "FALSE";
parameter LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE = "FALSE";
parameter [3:0] LINK_CTRL2_TARGET_LINK_SPEED = 4'h2;
parameter LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
parameter [14:0] LL_ACK_TIMEOUT = 15'h0000;
parameter LL_ACK_TIMEOUT_EN = "FALSE";
parameter LL_ACK_TIMEOUT_FUNC = 0;
parameter [14:0] LL_REPLAY_TIMEOUT = 15'h0000;
parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
parameter LL_REPLAY_TIMEOUT_FUNC = 0;
parameter [5:0] LTSSM_MAX_LINK_WIDTH = 6'h01;
parameter MPS_FORCE = "FALSE";
parameter [7:0] MSIX_BASE_PTR = 8'h9C;
parameter [7:0] MSIX_CAP_ID = 8'h11;
parameter [7:0] MSIX_CAP_NEXTPTR = 8'h00;
parameter MSIX_CAP_ON = "FALSE";
parameter MSIX_CAP_PBA_BIR = 0;
parameter [28:0] MSIX_CAP_PBA_OFFSET = 29'h00000050;
parameter MSIX_CAP_TABLE_BIR = 0;
parameter [28:0] MSIX_CAP_TABLE_OFFSET = 29'h00000040;
parameter [10:0] MSIX_CAP_TABLE_SIZE = 11'h000;
parameter [7:0] MSI_BASE_PTR = 8'h48;
parameter MSI_CAP_64_BIT_ADDR_CAPABLE = "TRUE";
parameter [7:0] MSI_CAP_ID = 8'h05;
parameter MSI_CAP_MULTIMSGCAP = 0;
parameter MSI_CAP_MULTIMSG_EXTENSION = 0;
parameter [7:0] MSI_CAP_NEXTPTR = 8'h60;
parameter MSI_CAP_ON = "FALSE";
parameter MSI_CAP_PER_VECTOR_MASKING_CAPABLE = "TRUE";
parameter N_FTS_COMCLK_GEN1 = 255;
parameter N_FTS_COMCLK_GEN2 = 255;
parameter N_FTS_GEN1 = 255;
parameter N_FTS_GEN2 = 255;
parameter [7:0] PCIE_BASE_PTR = 8'h60;
parameter [7:0] PCIE_CAP_CAPABILITY_ID = 8'h10;
parameter [3:0] PCIE_CAP_CAPABILITY_VERSION = 4'h2;
parameter [3:0] PCIE_CAP_DEVICE_PORT_TYPE = 4'h0;
parameter [7:0] PCIE_CAP_NEXTPTR = 8'h9C;
parameter PCIE_CAP_ON = "TRUE";
parameter PCIE_CAP_RSVD_15_14 = 0;
parameter PCIE_CAP_SLOT_IMPLEMENTED = "FALSE";
parameter PCIE_REVISION = 2;
parameter PL_AUTO_CONFIG = 0;
parameter PL_FAST_TRAIN = "FALSE";
parameter [14:0] PM_ASPML0S_TIMEOUT = 15'h0000;
parameter PM_ASPML0S_TIMEOUT_EN = "FALSE";
parameter PM_ASPML0S_TIMEOUT_FUNC = 0;
parameter PM_ASPM_FASTEXIT = "FALSE";
parameter [7:0] PM_BASE_PTR = 8'h40;
parameter PM_CAP_AUXCURRENT = 0;
parameter PM_CAP_D1SUPPORT = "TRUE";
parameter PM_CAP_D2SUPPORT = "TRUE";
parameter PM_CAP_DSI = "FALSE";
parameter [7:0] PM_CAP_ID = 8'h01;
parameter [7:0] PM_CAP_NEXTPTR = 8'h48;
parameter PM_CAP_ON = "TRUE";
parameter [4:0] PM_CAP_PMESUPPORT = 5'h0F;
parameter PM_CAP_PME_CLOCK = "FALSE";
parameter PM_CAP_RSVD_04 = 0;
parameter PM_CAP_VERSION = 3;
parameter PM_CSR_B2B3 = "FALSE";
parameter PM_CSR_BPCCEN = "FALSE";
parameter PM_CSR_NOSOFTRST = "TRUE";
parameter [7:0] PM_DATA0 = 8'h01;
parameter [7:0] PM_DATA1 = 8'h01;
parameter [7:0] PM_DATA2 = 8'h01;
parameter [7:0] PM_DATA3 = 8'h01;
parameter [7:0] PM_DATA4 = 8'h01;
parameter [7:0] PM_DATA5 = 8'h01;
parameter [7:0] PM_DATA6 = 8'h01;
parameter [7:0] PM_DATA7 = 8'h01;
parameter [1:0] PM_DATA_SCALE0 = 2'h1;
parameter [1:0] PM_DATA_SCALE1 = 2'h1;
parameter [1:0] PM_DATA_SCALE2 = 2'h1;
parameter [1:0] PM_DATA_SCALE3 = 2'h1;
parameter [1:0] PM_DATA_SCALE4 = 2'h1;
parameter [1:0] PM_DATA_SCALE5 = 2'h1;
parameter [1:0] PM_DATA_SCALE6 = 2'h1;
parameter [1:0] PM_DATA_SCALE7 = 2'h1;
parameter PM_MF = "FALSE";
parameter [11:0] RBAR_BASE_PTR = 12'h178;
parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR0 = 5'h00;
parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR1 = 5'h00;
parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR2 = 5'h00;
parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR3 = 5'h00;
parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR4 = 5'h00;
parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR5 = 5'h00;
parameter [15:0] RBAR_CAP_ID = 16'h0015;
parameter [2:0] RBAR_CAP_INDEX0 = 3'h0;
parameter [2:0] RBAR_CAP_INDEX1 = 3'h0;
parameter [2:0] RBAR_CAP_INDEX2 = 3'h0;
parameter [2:0] RBAR_CAP_INDEX3 = 3'h0;
parameter [2:0] RBAR_CAP_INDEX4 = 3'h0;
parameter [2:0] RBAR_CAP_INDEX5 = 3'h0;
parameter [11:0] RBAR_CAP_NEXTPTR = 12'h000;
parameter RBAR_CAP_ON = "FALSE";
parameter [31:0] RBAR_CAP_SUP0 = 32'h00000000;
parameter [31:0] RBAR_CAP_SUP1 = 32'h00000000;
parameter [31:0] RBAR_CAP_SUP2 = 32'h00000000;
parameter [31:0] RBAR_CAP_SUP3 = 32'h00000000;
parameter [31:0] RBAR_CAP_SUP4 = 32'h00000000;
parameter [31:0] RBAR_CAP_SUP5 = 32'h00000000;
parameter [3:0] RBAR_CAP_VERSION = 4'h1;
parameter [2:0] RBAR_NUM = 3'h1;
parameter RECRC_CHK = 0;
parameter RECRC_CHK_TRIM = "FALSE";
parameter ROOT_CAP_CRS_SW_VISIBILITY = "FALSE";
parameter [1:0] RP_AUTO_SPD = 2'h1;
parameter [4:0] RP_AUTO_SPD_LOOPCNT = 5'h1F;
parameter SELECT_DLL_IF = "FALSE";
parameter SIM_VERSION = "1.0";
parameter SLOT_CAP_ATT_BUTTON_PRESENT = "FALSE";
parameter SLOT_CAP_ATT_INDICATOR_PRESENT = "FALSE";
parameter SLOT_CAP_ELEC_INTERLOCK_PRESENT = "FALSE";
parameter SLOT_CAP_HOTPLUG_CAPABLE = "FALSE";
parameter SLOT_CAP_HOTPLUG_SURPRISE = "FALSE";
parameter SLOT_CAP_MRL_SENSOR_PRESENT = "FALSE";
parameter SLOT_CAP_NO_CMD_COMPLETED_SUPPORT = "FALSE";
parameter [12:0] SLOT_CAP_PHYSICAL_SLOT_NUM = 13'h0000;
parameter SLOT_CAP_POWER_CONTROLLER_PRESENT = "FALSE";
parameter SLOT_CAP_POWER_INDICATOR_PRESENT = "FALSE";
parameter SLOT_CAP_SLOT_POWER_LIMIT_SCALE = 0;
parameter [7:0] SLOT_CAP_SLOT_POWER_LIMIT_VALUE = 8'h00;
parameter SPARE_BIT0 = 0;
parameter SPARE_BIT1 = 0;
parameter SPARE_BIT2 = 0;
parameter SPARE_BIT3 = 0;
parameter SPARE_BIT4 = 0;
parameter SPARE_BIT5 = 0;
parameter SPARE_BIT6 = 0;
parameter SPARE_BIT7 = 0;
parameter SPARE_BIT8 = 0;
parameter [7:0] SPARE_BYTE0 = 8'h00;
parameter [7:0] SPARE_BYTE1 = 8'h00;
parameter [7:0] SPARE_BYTE2 = 8'h00;
parameter [7:0] SPARE_BYTE3 = 8'h00;
parameter [31:0] SPARE_WORD0 = 32'h00000000;
parameter [31:0] SPARE_WORD1 = 32'h00000000;
parameter [31:0] SPARE_WORD2 = 32'h00000000;
parameter [31:0] SPARE_WORD3 = 32'h00000000;
parameter SSL_MESSAGE_AUTO = "FALSE";
parameter TECRC_EP_INV = "FALSE";
parameter TL_RBYPASS = "FALSE";
parameter TL_RX_RAM_RADDR_LATENCY = 0;
parameter TL_RX_RAM_RDATA_LATENCY = 2;
parameter TL_RX_RAM_WRITE_LATENCY = 0;
parameter TL_TFC_DISABLE = "FALSE";
parameter TL_TX_CHECKS_DISABLE = "FALSE";
parameter TL_TX_RAM_RADDR_LATENCY = 0;
parameter TL_TX_RAM_RDATA_LATENCY = 2;
parameter TL_TX_RAM_WRITE_LATENCY = 0;
parameter TRN_DW = "FALSE";
parameter TRN_NP_FC = "FALSE";
parameter UPCONFIG_CAPABLE = "TRUE";
parameter UPSTREAM_FACING = "TRUE";
parameter UR_ATOMIC = "TRUE";
parameter UR_CFG1 = "TRUE";
parameter UR_INV_REQ = "TRUE";
parameter UR_PRS_RESPONSE = "TRUE";
parameter USER_CLK2_DIV2 = "FALSE";
parameter USER_CLK_FREQ = 3;
parameter USE_RID_PINS = "FALSE";
parameter VC0_CPL_INFINITE = "TRUE";
parameter [12:0] VC0_RX_RAM_LIMIT = 13'h03FF;
parameter VC0_TOTAL_CREDITS_CD = 127;
parameter VC0_TOTAL_CREDITS_CH = 31;
parameter VC0_TOTAL_CREDITS_NPD = 24;
parameter VC0_TOTAL_CREDITS_NPH = 12;
parameter VC0_TOTAL_CREDITS_PD = 288;
parameter VC0_TOTAL_CREDITS_PH = 32;
parameter VC0_TX_LASTPACKET = 31;
parameter [11:0] VC_BASE_PTR = 12'h10C;
parameter [15:0] VC_CAP_ID = 16'h0002;
parameter [11:0] VC_CAP_NEXTPTR = 12'h000;
parameter VC_CAP_ON = "FALSE";
parameter VC_CAP_REJECT_SNOOP_TRANSACTIONS = "FALSE";
parameter [3:0] VC_CAP_VERSION = 4'h1;
parameter [11:0] VSEC_BASE_PTR = 12'h128;
parameter [15:0] VSEC_CAP_HDR_ID = 16'h1234;
parameter [11:0] VSEC_CAP_HDR_LENGTH = 12'h018;
parameter [3:0] VSEC_CAP_HDR_REVISION = 4'h1;
parameter [15:0] VSEC_CAP_ID = 16'h000B;
parameter VSEC_CAP_IS_LINK_VISIBLE = "TRUE";
parameter [11:0] VSEC_CAP_NEXTPTR = 12'h140;
parameter VSEC_CAP_ON = "FALSE";
parameter [3:0] VSEC_CAP_VERSION = 4'h1;
endmodule
//#### END MODULE DEFINITION FOR: PCIE_2_1 ####

//#### BEGIN MODULE DEFINITION FOR :PCIE_3_0 ###
module PCIE_3_0 (
  CFGCURRENTSPEED,
  CFGDPASUBSTATECHANGE,
  CFGERRCOROUT,
  CFGERRFATALOUT,
  CFGERRNONFATALOUT,
  CFGEXTFUNCTIONNUMBER,
  CFGEXTREADRECEIVED,
  CFGEXTREGISTERNUMBER,
  CFGEXTWRITEBYTEENABLE,
  CFGEXTWRITEDATA,
  CFGEXTWRITERECEIVED,
  CFGFCCPLD,
  CFGFCCPLH,
  CFGFCNPD,
  CFGFCNPH,
  CFGFCPD,
  CFGFCPH,
  CFGFLRINPROCESS,
  CFGFUNCTIONPOWERSTATE,
  CFGFUNCTIONSTATUS,
  CFGHOTRESETOUT,
  CFGINPUTUPDATEDONE,
  CFGINTERRUPTAOUTPUT,
  CFGINTERRUPTBOUTPUT,
  CFGINTERRUPTCOUTPUT,
  CFGINTERRUPTDOUTPUT,
  CFGINTERRUPTMSIDATA,
  CFGINTERRUPTMSIENABLE,
  CFGINTERRUPTMSIFAIL,
  CFGINTERRUPTMSIMASKUPDATE,
  CFGINTERRUPTMSIMMENABLE,
  CFGINTERRUPTMSISENT,
  CFGINTERRUPTMSIVFENABLE,
  CFGINTERRUPTMSIXENABLE,
  CFGINTERRUPTMSIXFAIL,
  CFGINTERRUPTMSIXMASK,
  CFGINTERRUPTMSIXSENT,
  CFGINTERRUPTMSIXVFENABLE,
  CFGINTERRUPTMSIXVFMASK,
  CFGINTERRUPTSENT,
  CFGLINKPOWERSTATE,
  CFGLOCALERROR,
  CFGLTRENABLE,
  CFGLTSSMSTATE,
  CFGMAXPAYLOAD,
  CFGMAXREADREQ,
  CFGMCUPDATEDONE,
  CFGMGMTREADDATA,
  CFGMGMTREADWRITEDONE,
  CFGMSGRECEIVED,
  CFGMSGRECEIVEDDATA,
  CFGMSGRECEIVEDTYPE,
  CFGMSGTRANSMITDONE,
  CFGNEGOTIATEDWIDTH,
  CFGOBFFENABLE,
  CFGPERFUNCSTATUSDATA,
  CFGPERFUNCTIONUPDATEDONE,
  CFGPHYLINKDOWN,
  CFGPHYLINKSTATUS,
  CFGPLSTATUSCHANGE,
  CFGPOWERSTATECHANGEINTERRUPT,
  CFGRCBSTATUS,
  CFGTPHFUNCTIONNUM,
  CFGTPHREQUESTERENABLE,
  CFGTPHSTMODE,
  CFGTPHSTTADDRESS,
  CFGTPHSTTREADENABLE,
  CFGTPHSTTWRITEBYTEVALID,
  CFGTPHSTTWRITEDATA,
  CFGTPHSTTWRITEENABLE,
  CFGVFFLRINPROCESS,
  CFGVFPOWERSTATE,
  CFGVFSTATUS,
  CFGVFTPHREQUESTERENABLE,
  CFGVFTPHSTMODE,
  DBGDATAOUT,
  DRPDO,
  DRPRDY,
  MAXISCQTDATA,
  MAXISCQTKEEP,
  MAXISCQTLAST,
  MAXISCQTUSER,
  MAXISCQTVALID,
  MAXISRCTDATA,
  MAXISRCTKEEP,
  MAXISRCTLAST,
  MAXISRCTUSER,
  MAXISRCTVALID,
  MICOMPLETIONRAMREADADDRESSAL,
  MICOMPLETIONRAMREADADDRESSAU,
  MICOMPLETIONRAMREADADDRESSBL,
  MICOMPLETIONRAMREADADDRESSBU,
  MICOMPLETIONRAMREADENABLEL,
  MICOMPLETIONRAMREADENABLEU,
  MICOMPLETIONRAMWRITEADDRESSAL,
  MICOMPLETIONRAMWRITEADDRESSAU,
  MICOMPLETIONRAMWRITEADDRESSBL,
  MICOMPLETIONRAMWRITEADDRESSBU,
  MICOMPLETIONRAMWRITEDATAL,
  MICOMPLETIONRAMWRITEDATAU,
  MICOMPLETIONRAMWRITEENABLEL,
  MICOMPLETIONRAMWRITEENABLEU,
  MIREPLAYRAMADDRESS,
  MIREPLAYRAMREADENABLE,
  MIREPLAYRAMWRITEDATA,
  MIREPLAYRAMWRITEENABLE,
  MIREQUESTRAMREADADDRESSA,
  MIREQUESTRAMREADADDRESSB,
  MIREQUESTRAMREADENABLE,
  MIREQUESTRAMWRITEADDRESSA,
  MIREQUESTRAMWRITEADDRESSB,
  MIREQUESTRAMWRITEDATA,
  MIREQUESTRAMWRITEENABLE,
  PCIECQNPREQCOUNT,
  PCIERQSEQNUM,
  PCIERQSEQNUMVLD,
  PCIERQTAG,
  PCIERQTAGAV,
  PCIERQTAGVLD,
  PCIETFCNPDAV,
  PCIETFCNPHAV,
  PIPERX0EQCONTROL,
  PIPERX0EQLPLFFS,
  PIPERX0EQLPTXPRESET,
  PIPERX0EQPRESET,
  PIPERX0POLARITY,
  PIPERX1EQCONTROL,
  PIPERX1EQLPLFFS,
  PIPERX1EQLPTXPRESET,
  PIPERX1EQPRESET,
  PIPERX1POLARITY,
  PIPERX2EQCONTROL,
  PIPERX2EQLPLFFS,
  PIPERX2EQLPTXPRESET,
  PIPERX2EQPRESET,
  PIPERX2POLARITY,
  PIPERX3EQCONTROL,
  PIPERX3EQLPLFFS,
  PIPERX3EQLPTXPRESET,
  PIPERX3EQPRESET,
  PIPERX3POLARITY,
  PIPERX4EQCONTROL,
  PIPERX4EQLPLFFS,
  PIPERX4EQLPTXPRESET,
  PIPERX4EQPRESET,
  PIPERX4POLARITY,
  PIPERX5EQCONTROL,
  PIPERX5EQLPLFFS,
  PIPERX5EQLPTXPRESET,
  PIPERX5EQPRESET,
  PIPERX5POLARITY,
  PIPERX6EQCONTROL,
  PIPERX6EQLPLFFS,
  PIPERX6EQLPTXPRESET,
  PIPERX6EQPRESET,
  PIPERX6POLARITY,
  PIPERX7EQCONTROL,
  PIPERX7EQLPLFFS,
  PIPERX7EQLPTXPRESET,
  PIPERX7EQPRESET,
  PIPERX7POLARITY,
  PIPETX0CHARISK,
  PIPETX0COMPLIANCE,
  PIPETX0DATA,
  PIPETX0DATAVALID,
  PIPETX0ELECIDLE,
  PIPETX0EQCONTROL,
  PIPETX0EQDEEMPH,
  PIPETX0EQPRESET,
  PIPETX0POWERDOWN,
  PIPETX0STARTBLOCK,
  PIPETX0SYNCHEADER,
  PIPETX1CHARISK,
  PIPETX1COMPLIANCE,
  PIPETX1DATA,
  PIPETX1DATAVALID,
  PIPETX1ELECIDLE,
  PIPETX1EQCONTROL,
  PIPETX1EQDEEMPH,
  PIPETX1EQPRESET,
  PIPETX1POWERDOWN,
  PIPETX1STARTBLOCK,
  PIPETX1SYNCHEADER,
  PIPETX2CHARISK,
  PIPETX2COMPLIANCE,
  PIPETX2DATA,
  PIPETX2DATAVALID,
  PIPETX2ELECIDLE,
  PIPETX2EQCONTROL,
  PIPETX2EQDEEMPH,
  PIPETX2EQPRESET,
  PIPETX2POWERDOWN,
  PIPETX2STARTBLOCK,
  PIPETX2SYNCHEADER,
  PIPETX3CHARISK,
  PIPETX3COMPLIANCE,
  PIPETX3DATA,
  PIPETX3DATAVALID,
  PIPETX3ELECIDLE,
  PIPETX3EQCONTROL,
  PIPETX3EQDEEMPH,
  PIPETX3EQPRESET,
  PIPETX3POWERDOWN,
  PIPETX3STARTBLOCK,
  PIPETX3SYNCHEADER,
  PIPETX4CHARISK,
  PIPETX4COMPLIANCE,
  PIPETX4DATA,
  PIPETX4DATAVALID,
  PIPETX4ELECIDLE,
  PIPETX4EQCONTROL,
  PIPETX4EQDEEMPH,
  PIPETX4EQPRESET,
  PIPETX4POWERDOWN,
  PIPETX4STARTBLOCK,
  PIPETX4SYNCHEADER,
  PIPETX5CHARISK,
  PIPETX5COMPLIANCE,
  PIPETX5DATA,
  PIPETX5DATAVALID,
  PIPETX5ELECIDLE,
  PIPETX5EQCONTROL,
  PIPETX5EQDEEMPH,
  PIPETX5EQPRESET,
  PIPETX5POWERDOWN,
  PIPETX5STARTBLOCK,
  PIPETX5SYNCHEADER,
  PIPETX6CHARISK,
  PIPETX6COMPLIANCE,
  PIPETX6DATA,
  PIPETX6DATAVALID,
  PIPETX6ELECIDLE,
  PIPETX6EQCONTROL,
  PIPETX6EQDEEMPH,
  PIPETX6EQPRESET,
  PIPETX6POWERDOWN,
  PIPETX6STARTBLOCK,
  PIPETX6SYNCHEADER,
  PIPETX7CHARISK,
  PIPETX7COMPLIANCE,
  PIPETX7DATA,
  PIPETX7DATAVALID,
  PIPETX7ELECIDLE,
  PIPETX7EQCONTROL,
  PIPETX7EQDEEMPH,
  PIPETX7EQPRESET,
  PIPETX7POWERDOWN,
  PIPETX7STARTBLOCK,
  PIPETX7SYNCHEADER,
  PIPETXDEEMPH,
  PIPETXMARGIN,
  PIPETXRATE,
  PIPETXRCVRDET,
  PIPETXRESET,
  PIPETXSWING,
  PLEQINPROGRESS,
  PLEQPHASE,
  PLGEN3PCSRXSLIDE,
  SAXISCCTREADY,
  SAXISRQTREADY,

  CFGCONFIGSPACEENABLE,
  CFGDEVID,
  CFGDSBUSNUMBER,
  CFGDSDEVICENUMBER,
  CFGDSFUNCTIONNUMBER,
  CFGDSN,
  CFGDSPORTNUMBER,
  CFGERRCORIN,
  CFGERRUNCORIN,
  CFGEXTREADDATA,
  CFGEXTREADDATAVALID,
  CFGFCSEL,
  CFGFLRDONE,
  CFGHOTRESETIN,
  CFGINPUTUPDATEREQUEST,
  CFGINTERRUPTINT,
  CFGINTERRUPTMSIATTR,
  CFGINTERRUPTMSIFUNCTIONNUMBER,
  CFGINTERRUPTMSIINT,
  CFGINTERRUPTMSIPENDINGSTATUS,
  CFGINTERRUPTMSISELECT,
  CFGINTERRUPTMSITPHPRESENT,
  CFGINTERRUPTMSITPHSTTAG,
  CFGINTERRUPTMSITPHTYPE,
  CFGINTERRUPTMSIXADDRESS,
  CFGINTERRUPTMSIXDATA,
  CFGINTERRUPTMSIXINT,
  CFGINTERRUPTPENDING,
  CFGLINKTRAININGENABLE,
  CFGMCUPDATEREQUEST,
  CFGMGMTADDR,
  CFGMGMTBYTEENABLE,
  CFGMGMTREAD,
  CFGMGMTTYPE1CFGREGACCESS,
  CFGMGMTWRITE,
  CFGMGMTWRITEDATA,
  CFGMSGTRANSMIT,
  CFGMSGTRANSMITDATA,
  CFGMSGTRANSMITTYPE,
  CFGPERFUNCSTATUSCONTROL,
  CFGPERFUNCTIONNUMBER,
  CFGPERFUNCTIONOUTPUTREQUEST,
  CFGPOWERSTATECHANGEACK,
  CFGREQPMTRANSITIONL23READY,
  CFGREVID,
  CFGSUBSYSID,
  CFGSUBSYSVENDID,
  CFGTPHSTTREADDATA,
  CFGTPHSTTREADDATAVALID,
  CFGVENDID,
  CFGVFFLRDONE,
  CORECLK,
  CORECLKMICOMPLETIONRAML,
  CORECLKMICOMPLETIONRAMU,
  CORECLKMIREPLAYRAM,
  CORECLKMIREQUESTRAM,
  DRPADDR,
  DRPCLK,
  DRPDI,
  DRPEN,
  DRPWE,
  MAXISCQTREADY,
  MAXISRCTREADY,
  MGMTRESETN,
  MGMTSTICKYRESETN,
  MICOMPLETIONRAMREADDATA,
  MIREPLAYRAMREADDATA,
  MIREQUESTRAMREADDATA,
  PCIECQNPREQ,
  PIPECLK,
  PIPEEQFS,
  PIPEEQLF,
  PIPERESETN,
  PIPERX0CHARISK,
  PIPERX0DATA,
  PIPERX0DATAVALID,
  PIPERX0ELECIDLE,
  PIPERX0EQDONE,
  PIPERX0EQLPADAPTDONE,
  PIPERX0EQLPLFFSSEL,
  PIPERX0EQLPNEWTXCOEFFORPRESET,
  PIPERX0PHYSTATUS,
  PIPERX0STARTBLOCK,
  PIPERX0STATUS,
  PIPERX0SYNCHEADER,
  PIPERX0VALID,
  PIPERX1CHARISK,
  PIPERX1DATA,
  PIPERX1DATAVALID,
  PIPERX1ELECIDLE,
  PIPERX1EQDONE,
  PIPERX1EQLPADAPTDONE,
  PIPERX1EQLPLFFSSEL,
  PIPERX1EQLPNEWTXCOEFFORPRESET,
  PIPERX1PHYSTATUS,
  PIPERX1STARTBLOCK,
  PIPERX1STATUS,
  PIPERX1SYNCHEADER,
  PIPERX1VALID,
  PIPERX2CHARISK,
  PIPERX2DATA,
  PIPERX2DATAVALID,
  PIPERX2ELECIDLE,
  PIPERX2EQDONE,
  PIPERX2EQLPADAPTDONE,
  PIPERX2EQLPLFFSSEL,
  PIPERX2EQLPNEWTXCOEFFORPRESET,
  PIPERX2PHYSTATUS,
  PIPERX2STARTBLOCK,
  PIPERX2STATUS,
  PIPERX2SYNCHEADER,
  PIPERX2VALID,
  PIPERX3CHARISK,
  PIPERX3DATA,
  PIPERX3DATAVALID,
  PIPERX3ELECIDLE,
  PIPERX3EQDONE,
  PIPERX3EQLPADAPTDONE,
  PIPERX3EQLPLFFSSEL,
  PIPERX3EQLPNEWTXCOEFFORPRESET,
  PIPERX3PHYSTATUS,
  PIPERX3STARTBLOCK,
  PIPERX3STATUS,
  PIPERX3SYNCHEADER,
  PIPERX3VALID,
  PIPERX4CHARISK,
  PIPERX4DATA,
  PIPERX4DATAVALID,
  PIPERX4ELECIDLE,
  PIPERX4EQDONE,
  PIPERX4EQLPADAPTDONE,
  PIPERX4EQLPLFFSSEL,
  PIPERX4EQLPNEWTXCOEFFORPRESET,
  PIPERX4PHYSTATUS,
  PIPERX4STARTBLOCK,
  PIPERX4STATUS,
  PIPERX4SYNCHEADER,
  PIPERX4VALID,
  PIPERX5CHARISK,
  PIPERX5DATA,
  PIPERX5DATAVALID,
  PIPERX5ELECIDLE,
  PIPERX5EQDONE,
  PIPERX5EQLPADAPTDONE,
  PIPERX5EQLPLFFSSEL,
  PIPERX5EQLPNEWTXCOEFFORPRESET,
  PIPERX5PHYSTATUS,
  PIPERX5STARTBLOCK,
  PIPERX5STATUS,
  PIPERX5SYNCHEADER,
  PIPERX5VALID,
  PIPERX6CHARISK,
  PIPERX6DATA,
  PIPERX6DATAVALID,
  PIPERX6ELECIDLE,
  PIPERX6EQDONE,
  PIPERX6EQLPADAPTDONE,
  PIPERX6EQLPLFFSSEL,
  PIPERX6EQLPNEWTXCOEFFORPRESET,
  PIPERX6PHYSTATUS,
  PIPERX6STARTBLOCK,
  PIPERX6STATUS,
  PIPERX6SYNCHEADER,
  PIPERX6VALID,
  PIPERX7CHARISK,
  PIPERX7DATA,
  PIPERX7DATAVALID,
  PIPERX7ELECIDLE,
  PIPERX7EQDONE,
  PIPERX7EQLPADAPTDONE,
  PIPERX7EQLPLFFSSEL,
  PIPERX7EQLPNEWTXCOEFFORPRESET,
  PIPERX7PHYSTATUS,
  PIPERX7STARTBLOCK,
  PIPERX7STATUS,
  PIPERX7SYNCHEADER,
  PIPERX7VALID,
  PIPETX0EQCOEFF,
  PIPETX0EQDONE,
  PIPETX1EQCOEFF,
  PIPETX1EQDONE,
  PIPETX2EQCOEFF,
  PIPETX2EQDONE,
  PIPETX3EQCOEFF,
  PIPETX3EQDONE,
  PIPETX4EQCOEFF,
  PIPETX4EQDONE,
  PIPETX5EQCOEFF,
  PIPETX5EQDONE,
  PIPETX6EQCOEFF,
  PIPETX6EQDONE,
  PIPETX7EQCOEFF,
  PIPETX7EQDONE,
  PLDISABLESCRAMBLER,
  PLEQRESETEIEOSCOUNT,
  PLGEN3PCSDISABLE,
  PLGEN3PCSRXSYNCDONE,
  RECCLK,
  RESETN,
  SAXISCCTDATA,
  SAXISCCTKEEP,
  SAXISCCTLAST,
  SAXISCCTUSER,
  SAXISCCTVALID,
  SAXISRQTDATA,
  SAXISRQTKEEP,
  SAXISRQTLAST,
  SAXISRQTUSER,
  SAXISRQTVALID,
  USERCLK
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CFGCONFIGSPACEENABLE ;
input CFGERRCORIN ;
input CFGERRUNCORIN ;
input CFGEXTREADDATAVALID ;
input CFGHOTRESETIN ;
input CFGINPUTUPDATEREQUEST ;
input CFGINTERRUPTMSITPHPRESENT ;
input CFGINTERRUPTMSIXINT ;
input CFGLINKTRAININGENABLE ;
input CFGMCUPDATEREQUEST ;
input CFGMGMTREAD ;
input CFGMGMTTYPE1CFGREGACCESS ;
input CFGMGMTWRITE ;
input CFGMSGTRANSMIT ;
input CFGPERFUNCTIONOUTPUTREQUEST ;
input CFGPOWERSTATECHANGEACK ;
input CFGREQPMTRANSITIONL23READY ;
input CFGTPHSTTREADDATAVALID ;
input CORECLK ;
input CORECLKMICOMPLETIONRAML ;
input CORECLKMICOMPLETIONRAMU ;
input CORECLKMIREPLAYRAM ;
input CORECLKMIREQUESTRAM ;
input DRPCLK ;
input DRPEN ;
input DRPWE ;
input MGMTRESETN ;
input MGMTSTICKYRESETN ;
input PCIECQNPREQ ;
input PIPECLK ;
input PIPERESETN ;
input PIPERX0DATAVALID ;
input PIPERX0ELECIDLE ;
input PIPERX0EQDONE ;
input PIPERX0EQLPADAPTDONE ;
input PIPERX0EQLPLFFSSEL ;
input PIPERX0PHYSTATUS ;
input PIPERX0STARTBLOCK ;
input PIPERX0VALID ;
input PIPERX1DATAVALID ;
input PIPERX1ELECIDLE ;
input PIPERX1EQDONE ;
input PIPERX1EQLPADAPTDONE ;
input PIPERX1EQLPLFFSSEL ;
input PIPERX1PHYSTATUS ;
input PIPERX1STARTBLOCK ;
input PIPERX1VALID ;
input PIPERX2DATAVALID ;
input PIPERX2ELECIDLE ;
input PIPERX2EQDONE ;
input PIPERX2EQLPADAPTDONE ;
input PIPERX2EQLPLFFSSEL ;
input PIPERX2PHYSTATUS ;
input PIPERX2STARTBLOCK ;
input PIPERX2VALID ;
input PIPERX3DATAVALID ;
input PIPERX3ELECIDLE ;
input PIPERX3EQDONE ;
input PIPERX3EQLPADAPTDONE ;
input PIPERX3EQLPLFFSSEL ;
input PIPERX3PHYSTATUS ;
input PIPERX3STARTBLOCK ;
input PIPERX3VALID ;
input PIPERX4DATAVALID ;
input PIPERX4ELECIDLE ;
input PIPERX4EQDONE ;
input PIPERX4EQLPADAPTDONE ;
input PIPERX4EQLPLFFSSEL ;
input PIPERX4PHYSTATUS ;
input PIPERX4STARTBLOCK ;
input PIPERX4VALID ;
input PIPERX5DATAVALID ;
input PIPERX5ELECIDLE ;
input PIPERX5EQDONE ;
input PIPERX5EQLPADAPTDONE ;
input PIPERX5EQLPLFFSSEL ;
input PIPERX5PHYSTATUS ;
input PIPERX5STARTBLOCK ;
input PIPERX5VALID ;
input PIPERX6DATAVALID ;
input PIPERX6ELECIDLE ;
input PIPERX6EQDONE ;
input PIPERX6EQLPADAPTDONE ;
input PIPERX6EQLPLFFSSEL ;
input PIPERX6PHYSTATUS ;
input PIPERX6STARTBLOCK ;
input PIPERX6VALID ;
input PIPERX7DATAVALID ;
input PIPERX7ELECIDLE ;
input PIPERX7EQDONE ;
input PIPERX7EQLPADAPTDONE ;
input PIPERX7EQLPLFFSSEL ;
input PIPERX7PHYSTATUS ;
input PIPERX7STARTBLOCK ;
input PIPERX7VALID ;
input PIPETX0EQDONE ;
input PIPETX1EQDONE ;
input PIPETX2EQDONE ;
input PIPETX3EQDONE ;
input PIPETX4EQDONE ;
input PIPETX5EQDONE ;
input PIPETX6EQDONE ;
input PIPETX7EQDONE ;
input PLDISABLESCRAMBLER ;
input PLEQRESETEIEOSCOUNT ;
input PLGEN3PCSDISABLE ;
input RECCLK ;
input RESETN ;
input SAXISCCTLAST ;
input SAXISCCTVALID ;
input SAXISRQTLAST ;
input SAXISRQTVALID ;
input USERCLK ;
input [10:0] DRPADDR ;
input [143:0] MICOMPLETIONRAMREADDATA ;
input [143:0] MIREPLAYRAMREADDATA ;
input [143:0] MIREQUESTRAMREADDATA ;
input [15:0] CFGDEVID ;
input [15:0] CFGSUBSYSID ;
input [15:0] CFGSUBSYSVENDID ;
input [15:0] CFGVENDID ;
input [15:0] DRPDI ;
input [17:0] PIPERX0EQLPNEWTXCOEFFORPRESET ;
input [17:0] PIPERX1EQLPNEWTXCOEFFORPRESET ;
input [17:0] PIPERX2EQLPNEWTXCOEFFORPRESET ;
input [17:0] PIPERX3EQLPNEWTXCOEFFORPRESET ;
input [17:0] PIPERX4EQLPNEWTXCOEFFORPRESET ;
input [17:0] PIPERX5EQLPNEWTXCOEFFORPRESET ;
input [17:0] PIPERX6EQLPNEWTXCOEFFORPRESET ;
input [17:0] PIPERX7EQLPNEWTXCOEFFORPRESET ;
input [17:0] PIPETX0EQCOEFF ;
input [17:0] PIPETX1EQCOEFF ;
input [17:0] PIPETX2EQCOEFF ;
input [17:0] PIPETX3EQCOEFF ;
input [17:0] PIPETX4EQCOEFF ;
input [17:0] PIPETX5EQCOEFF ;
input [17:0] PIPETX6EQCOEFF ;
input [17:0] PIPETX7EQCOEFF ;
input [18:0] CFGMGMTADDR ;
input [1:0] CFGFLRDONE ;
input [1:0] CFGINTERRUPTMSITPHTYPE ;
input [1:0] CFGINTERRUPTPENDING ;
input [1:0] PIPERX0CHARISK ;
input [1:0] PIPERX0SYNCHEADER ;
input [1:0] PIPERX1CHARISK ;
input [1:0] PIPERX1SYNCHEADER ;
input [1:0] PIPERX2CHARISK ;
input [1:0] PIPERX2SYNCHEADER ;
input [1:0] PIPERX3CHARISK ;
input [1:0] PIPERX3SYNCHEADER ;
input [1:0] PIPERX4CHARISK ;
input [1:0] PIPERX4SYNCHEADER ;
input [1:0] PIPERX5CHARISK ;
input [1:0] PIPERX5SYNCHEADER ;
input [1:0] PIPERX6CHARISK ;
input [1:0] PIPERX6SYNCHEADER ;
input [1:0] PIPERX7CHARISK ;
input [1:0] PIPERX7SYNCHEADER ;
input [21:0] MAXISCQTREADY ;
input [21:0] MAXISRCTREADY ;
input [255:0] SAXISCCTDATA ;
input [255:0] SAXISRQTDATA ;
input [2:0] CFGDSFUNCTIONNUMBER ;
input [2:0] CFGFCSEL ;
input [2:0] CFGINTERRUPTMSIATTR ;
input [2:0] CFGINTERRUPTMSIFUNCTIONNUMBER ;
input [2:0] CFGMSGTRANSMITTYPE ;
input [2:0] CFGPERFUNCSTATUSCONTROL ;
input [2:0] CFGPERFUNCTIONNUMBER ;
input [2:0] PIPERX0STATUS ;
input [2:0] PIPERX1STATUS ;
input [2:0] PIPERX2STATUS ;
input [2:0] PIPERX3STATUS ;
input [2:0] PIPERX4STATUS ;
input [2:0] PIPERX5STATUS ;
input [2:0] PIPERX6STATUS ;
input [2:0] PIPERX7STATUS ;
input [31:0] CFGEXTREADDATA ;
input [31:0] CFGINTERRUPTMSIINT ;
input [31:0] CFGINTERRUPTMSIXDATA ;
input [31:0] CFGMGMTWRITEDATA ;
input [31:0] CFGMSGTRANSMITDATA ;
input [31:0] CFGTPHSTTREADDATA ;
input [31:0] PIPERX0DATA ;
input [31:0] PIPERX1DATA ;
input [31:0] PIPERX2DATA ;
input [31:0] PIPERX3DATA ;
input [31:0] PIPERX4DATA ;
input [31:0] PIPERX5DATA ;
input [31:0] PIPERX6DATA ;
input [31:0] PIPERX7DATA ;
input [32:0] SAXISCCTUSER ;
input [3:0] CFGINTERRUPTINT ;
input [3:0] CFGINTERRUPTMSISELECT ;
input [3:0] CFGMGMTBYTEENABLE ;
input [4:0] CFGDSDEVICENUMBER ;
input [59:0] SAXISRQTUSER ;
input [5:0] CFGVFFLRDONE ;
input [5:0] PIPEEQFS ;
input [5:0] PIPEEQLF ;
input [63:0] CFGDSN ;
input [63:0] CFGINTERRUPTMSIPENDINGSTATUS ;
input [63:0] CFGINTERRUPTMSIXADDRESS ;
input [7:0] CFGDSBUSNUMBER ;
input [7:0] CFGDSPORTNUMBER ;
input [7:0] CFGREVID ;
input [7:0] PLGEN3PCSRXSYNCDONE ;
input [7:0] SAXISCCTKEEP ;
input [7:0] SAXISRQTKEEP ;
input [8:0] CFGINTERRUPTMSITPHSTTAG ;
output CFGERRCOROUT ;
output CFGERRFATALOUT ;
output CFGERRNONFATALOUT ;
output CFGEXTREADRECEIVED ;
output CFGEXTWRITERECEIVED ;
output CFGHOTRESETOUT ;
output CFGINPUTUPDATEDONE ;
output CFGINTERRUPTAOUTPUT ;
output CFGINTERRUPTBOUTPUT ;
output CFGINTERRUPTCOUTPUT ;
output CFGINTERRUPTDOUTPUT ;
output CFGINTERRUPTMSIFAIL ;
output CFGINTERRUPTMSIMASKUPDATE ;
output CFGINTERRUPTMSISENT ;
output CFGINTERRUPTMSIXFAIL ;
output CFGINTERRUPTMSIXSENT ;
output CFGINTERRUPTSENT ;
output CFGLOCALERROR ;
output CFGLTRENABLE ;
output CFGMCUPDATEDONE ;
output CFGMGMTREADWRITEDONE ;
output CFGMSGRECEIVED ;
output CFGMSGTRANSMITDONE ;
output CFGPERFUNCTIONUPDATEDONE ;
output CFGPHYLINKDOWN ;
output CFGPLSTATUSCHANGE ;
output CFGPOWERSTATECHANGEINTERRUPT ;
output CFGTPHSTTREADENABLE ;
output CFGTPHSTTWRITEENABLE ;
output DRPRDY ;
output MAXISCQTLAST ;
output MAXISCQTVALID ;
output MAXISRCTLAST ;
output MAXISRCTVALID ;
output PCIERQSEQNUMVLD ;
output PCIERQTAGVLD ;
output PIPERX0POLARITY ;
output PIPERX1POLARITY ;
output PIPERX2POLARITY ;
output PIPERX3POLARITY ;
output PIPERX4POLARITY ;
output PIPERX5POLARITY ;
output PIPERX6POLARITY ;
output PIPERX7POLARITY ;
output PIPETX0COMPLIANCE ;
output PIPETX0DATAVALID ;
output PIPETX0ELECIDLE ;
output PIPETX0STARTBLOCK ;
output PIPETX1COMPLIANCE ;
output PIPETX1DATAVALID ;
output PIPETX1ELECIDLE ;
output PIPETX1STARTBLOCK ;
output PIPETX2COMPLIANCE ;
output PIPETX2DATAVALID ;
output PIPETX2ELECIDLE ;
output PIPETX2STARTBLOCK ;
output PIPETX3COMPLIANCE ;
output PIPETX3DATAVALID ;
output PIPETX3ELECIDLE ;
output PIPETX3STARTBLOCK ;
output PIPETX4COMPLIANCE ;
output PIPETX4DATAVALID ;
output PIPETX4ELECIDLE ;
output PIPETX4STARTBLOCK ;
output PIPETX5COMPLIANCE ;
output PIPETX5DATAVALID ;
output PIPETX5ELECIDLE ;
output PIPETX5STARTBLOCK ;
output PIPETX6COMPLIANCE ;
output PIPETX6DATAVALID ;
output PIPETX6ELECIDLE ;
output PIPETX6STARTBLOCK ;
output PIPETX7COMPLIANCE ;
output PIPETX7DATAVALID ;
output PIPETX7ELECIDLE ;
output PIPETX7STARTBLOCK ;
output PIPETXDEEMPH ;
output PIPETXRCVRDET ;
output PIPETXRESET ;
output PIPETXSWING ;
output PLEQINPROGRESS ;
output [11:0] CFGFCCPLD ;
output [11:0] CFGFCNPD ;
output [11:0] CFGFCPD ;
output [11:0] CFGVFSTATUS ;
output [143:0] MIREPLAYRAMWRITEDATA ;
output [143:0] MIREQUESTRAMWRITEDATA ;
output [15:0] CFGPERFUNCSTATUSDATA ;
output [15:0] DBGDATAOUT ;
output [15:0] DRPDO ;
output [17:0] CFGVFPOWERSTATE ;
output [17:0] CFGVFTPHSTMODE ;
output [1:0] CFGDPASUBSTATECHANGE ;
output [1:0] CFGFLRINPROCESS ;
output [1:0] CFGINTERRUPTMSIENABLE ;
output [1:0] CFGINTERRUPTMSIXENABLE ;
output [1:0] CFGINTERRUPTMSIXMASK ;
output [1:0] CFGLINKPOWERSTATE ;
output [1:0] CFGOBFFENABLE ;
output [1:0] CFGPHYLINKSTATUS ;
output [1:0] CFGRCBSTATUS ;
output [1:0] CFGTPHREQUESTERENABLE ;
output [1:0] MIREPLAYRAMREADENABLE ;
output [1:0] MIREPLAYRAMWRITEENABLE ;
output [1:0] PCIERQTAGAV ;
output [1:0] PCIETFCNPDAV ;
output [1:0] PCIETFCNPHAV ;
output [1:0] PIPERX0EQCONTROL ;
output [1:0] PIPERX1EQCONTROL ;
output [1:0] PIPERX2EQCONTROL ;
output [1:0] PIPERX3EQCONTROL ;
output [1:0] PIPERX4EQCONTROL ;
output [1:0] PIPERX5EQCONTROL ;
output [1:0] PIPERX6EQCONTROL ;
output [1:0] PIPERX7EQCONTROL ;
output [1:0] PIPETX0CHARISK ;
output [1:0] PIPETX0EQCONTROL ;
output [1:0] PIPETX0POWERDOWN ;
output [1:0] PIPETX0SYNCHEADER ;
output [1:0] PIPETX1CHARISK ;
output [1:0] PIPETX1EQCONTROL ;
output [1:0] PIPETX1POWERDOWN ;
output [1:0] PIPETX1SYNCHEADER ;
output [1:0] PIPETX2CHARISK ;
output [1:0] PIPETX2EQCONTROL ;
output [1:0] PIPETX2POWERDOWN ;
output [1:0] PIPETX2SYNCHEADER ;
output [1:0] PIPETX3CHARISK ;
output [1:0] PIPETX3EQCONTROL ;
output [1:0] PIPETX3POWERDOWN ;
output [1:0] PIPETX3SYNCHEADER ;
output [1:0] PIPETX4CHARISK ;
output [1:0] PIPETX4EQCONTROL ;
output [1:0] PIPETX4POWERDOWN ;
output [1:0] PIPETX4SYNCHEADER ;
output [1:0] PIPETX5CHARISK ;
output [1:0] PIPETX5EQCONTROL ;
output [1:0] PIPETX5POWERDOWN ;
output [1:0] PIPETX5SYNCHEADER ;
output [1:0] PIPETX6CHARISK ;
output [1:0] PIPETX6EQCONTROL ;
output [1:0] PIPETX6POWERDOWN ;
output [1:0] PIPETX6SYNCHEADER ;
output [1:0] PIPETX7CHARISK ;
output [1:0] PIPETX7EQCONTROL ;
output [1:0] PIPETX7POWERDOWN ;
output [1:0] PIPETX7SYNCHEADER ;
output [1:0] PIPETXRATE ;
output [1:0] PLEQPHASE ;
output [255:0] MAXISCQTDATA ;
output [255:0] MAXISRCTDATA ;
output [2:0] CFGCURRENTSPEED ;
output [2:0] CFGMAXPAYLOAD ;
output [2:0] CFGMAXREADREQ ;
output [2:0] CFGTPHFUNCTIONNUM ;
output [2:0] PIPERX0EQPRESET ;
output [2:0] PIPERX1EQPRESET ;
output [2:0] PIPERX2EQPRESET ;
output [2:0] PIPERX3EQPRESET ;
output [2:0] PIPERX4EQPRESET ;
output [2:0] PIPERX5EQPRESET ;
output [2:0] PIPERX6EQPRESET ;
output [2:0] PIPERX7EQPRESET ;
output [2:0] PIPETXMARGIN ;
output [31:0] CFGEXTWRITEDATA ;
output [31:0] CFGINTERRUPTMSIDATA ;
output [31:0] CFGMGMTREADDATA ;
output [31:0] CFGTPHSTTWRITEDATA ;
output [31:0] PIPETX0DATA ;
output [31:0] PIPETX1DATA ;
output [31:0] PIPETX2DATA ;
output [31:0] PIPETX3DATA ;
output [31:0] PIPETX4DATA ;
output [31:0] PIPETX5DATA ;
output [31:0] PIPETX6DATA ;
output [31:0] PIPETX7DATA ;
output [3:0] CFGEXTWRITEBYTEENABLE ;
output [3:0] CFGNEGOTIATEDWIDTH ;
output [3:0] CFGTPHSTTWRITEBYTEVALID ;
output [3:0] MICOMPLETIONRAMREADENABLEL ;
output [3:0] MICOMPLETIONRAMREADENABLEU ;
output [3:0] MICOMPLETIONRAMWRITEENABLEL ;
output [3:0] MICOMPLETIONRAMWRITEENABLEU ;
output [3:0] MIREQUESTRAMREADENABLE ;
output [3:0] MIREQUESTRAMWRITEENABLE ;
output [3:0] PCIERQSEQNUM ;
output [3:0] PIPERX0EQLPTXPRESET ;
output [3:0] PIPERX1EQLPTXPRESET ;
output [3:0] PIPERX2EQLPTXPRESET ;
output [3:0] PIPERX3EQLPTXPRESET ;
output [3:0] PIPERX4EQLPTXPRESET ;
output [3:0] PIPERX5EQLPTXPRESET ;
output [3:0] PIPERX6EQLPTXPRESET ;
output [3:0] PIPERX7EQLPTXPRESET ;
output [3:0] PIPETX0EQPRESET ;
output [3:0] PIPETX1EQPRESET ;
output [3:0] PIPETX2EQPRESET ;
output [3:0] PIPETX3EQPRESET ;
output [3:0] PIPETX4EQPRESET ;
output [3:0] PIPETX5EQPRESET ;
output [3:0] PIPETX6EQPRESET ;
output [3:0] PIPETX7EQPRESET ;
output [3:0] SAXISCCTREADY ;
output [3:0] SAXISRQTREADY ;
output [4:0] CFGMSGRECEIVEDTYPE ;
output [4:0] CFGTPHSTTADDRESS ;
output [5:0] CFGFUNCTIONPOWERSTATE ;
output [5:0] CFGINTERRUPTMSIMMENABLE ;
output [5:0] CFGINTERRUPTMSIVFENABLE ;
output [5:0] CFGINTERRUPTMSIXVFENABLE ;
output [5:0] CFGINTERRUPTMSIXVFMASK ;
output [5:0] CFGLTSSMSTATE ;
output [5:0] CFGTPHSTMODE ;
output [5:0] CFGVFFLRINPROCESS ;
output [5:0] CFGVFTPHREQUESTERENABLE ;
output [5:0] PCIECQNPREQCOUNT ;
output [5:0] PCIERQTAG ;
output [5:0] PIPERX0EQLPLFFS ;
output [5:0] PIPERX1EQLPLFFS ;
output [5:0] PIPERX2EQLPLFFS ;
output [5:0] PIPERX3EQLPLFFS ;
output [5:0] PIPERX4EQLPLFFS ;
output [5:0] PIPERX5EQLPLFFS ;
output [5:0] PIPERX6EQLPLFFS ;
output [5:0] PIPERX7EQLPLFFS ;
output [5:0] PIPETX0EQDEEMPH ;
output [5:0] PIPETX1EQDEEMPH ;
output [5:0] PIPETX2EQDEEMPH ;
output [5:0] PIPETX3EQDEEMPH ;
output [5:0] PIPETX4EQDEEMPH ;
output [5:0] PIPETX5EQDEEMPH ;
output [5:0] PIPETX6EQDEEMPH ;
output [5:0] PIPETX7EQDEEMPH ;
output [71:0] MICOMPLETIONRAMWRITEDATAL ;
output [71:0] MICOMPLETIONRAMWRITEDATAU ;
output [74:0] MAXISRCTUSER ;
output [7:0] CFGEXTFUNCTIONNUMBER ;
output [7:0] CFGFCCPLH ;
output [7:0] CFGFCNPH ;
output [7:0] CFGFCPH ;
output [7:0] CFGFUNCTIONSTATUS ;
output [7:0] CFGMSGRECEIVEDDATA ;
output [7:0] MAXISCQTKEEP ;
output [7:0] MAXISRCTKEEP ;
output [7:0] PLGEN3PCSRXSLIDE ;
output [84:0] MAXISCQTUSER ;
output [8:0] MIREPLAYRAMADDRESS ;
output [8:0] MIREQUESTRAMREADADDRESSA ;
output [8:0] MIREQUESTRAMREADADDRESSB ;
output [8:0] MIREQUESTRAMWRITEADDRESSA ;
output [8:0] MIREQUESTRAMWRITEADDRESSB ;
output [9:0] CFGEXTREGISTERNUMBER ;
output [9:0] MICOMPLETIONRAMREADADDRESSAL ;
output [9:0] MICOMPLETIONRAMREADADDRESSAU ;
output [9:0] MICOMPLETIONRAMREADADDRESSBL ;
output [9:0] MICOMPLETIONRAMREADADDRESSBU ;
output [9:0] MICOMPLETIONRAMWRITEADDRESSAL ;
output [9:0] MICOMPLETIONRAMWRITEADDRESSAU ;
output [9:0] MICOMPLETIONRAMWRITEADDRESSBL ;
output [9:0] MICOMPLETIONRAMWRITEADDRESSBU ;
parameter ARI_CAP_ENABLE = "FALSE";
parameter AXISTEN_IF_CC_ALIGNMENT_MODE = "FALSE";
parameter AXISTEN_IF_CC_PARITY_CHK = "TRUE";
parameter AXISTEN_IF_CQ_ALIGNMENT_MODE = "FALSE";
parameter AXISTEN_IF_ENABLE_CLIENT_TAG = "FALSE";
parameter [17:0] AXISTEN_IF_ENABLE_MSG_ROUTE = 18'h00000;
parameter AXISTEN_IF_ENABLE_RX_MSG_INTFC = "FALSE";
parameter AXISTEN_IF_RC_ALIGNMENT_MODE = "FALSE";
parameter AXISTEN_IF_RC_STRADDLE = "FALSE";
parameter AXISTEN_IF_RQ_ALIGNMENT_MODE = "FALSE";
parameter AXISTEN_IF_RQ_PARITY_CHK = "TRUE";
parameter [1:0] AXISTEN_IF_WIDTH = 2'h2;
parameter CRM_CORE_CLK_FREQ_500 = "TRUE";
parameter [1:0] CRM_USER_CLK_FREQ = 2'h2;
parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
parameter [1:0] GEN3_PCS_AUTO_REALIGN = 2'h1;
parameter GEN3_PCS_RX_ELECIDLE_INTERNAL = "TRUE";
parameter [8:0] LL_ACK_TIMEOUT = 9'h000;
parameter LL_ACK_TIMEOUT_EN = "FALSE";
parameter LL_ACK_TIMEOUT_FUNC = 0;
parameter [15:0] LL_CPL_FC_UPDATE_TIMER = 16'h0000;
parameter LL_CPL_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
parameter [15:0] LL_FC_UPDATE_TIMER = 16'h0000;
parameter LL_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
parameter [15:0] LL_NP_FC_UPDATE_TIMER = 16'h0000;
parameter LL_NP_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
parameter [15:0] LL_P_FC_UPDATE_TIMER = 16'h0000;
parameter LL_P_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
parameter [8:0] LL_REPLAY_TIMEOUT = 9'h000;
parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
parameter LL_REPLAY_TIMEOUT_FUNC = 0;
parameter [9:0] LTR_TX_MESSAGE_MINIMUM_INTERVAL = 10'h0FA;
parameter LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE = "FALSE";
parameter LTR_TX_MESSAGE_ON_LTR_ENABLE = "FALSE";
parameter PF0_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
parameter PF0_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
parameter [11:0] PF0_AER_CAP_NEXTPTR = 12'h000;
parameter [11:0] PF0_ARI_CAP_NEXTPTR = 12'h000;
parameter [7:0] PF0_ARI_CAP_NEXT_FUNC = 8'h00;
parameter [3:0] PF0_ARI_CAP_VER = 4'h1;
parameter [4:0] PF0_BAR0_APERTURE_SIZE = 5'h03;
parameter [2:0] PF0_BAR0_CONTROL = 3'h4;
parameter [4:0] PF0_BAR1_APERTURE_SIZE = 5'h00;
parameter [2:0] PF0_BAR1_CONTROL = 3'h0;
parameter [4:0] PF0_BAR2_APERTURE_SIZE = 5'h03;
parameter [2:0] PF0_BAR2_CONTROL = 3'h4;
parameter [4:0] PF0_BAR3_APERTURE_SIZE = 5'h03;
parameter [2:0] PF0_BAR3_CONTROL = 3'h0;
parameter [4:0] PF0_BAR4_APERTURE_SIZE = 5'h03;
parameter [2:0] PF0_BAR4_CONTROL = 3'h4;
parameter [4:0] PF0_BAR5_APERTURE_SIZE = 5'h03;
parameter [2:0] PF0_BAR5_CONTROL = 3'h0;
parameter [7:0] PF0_BIST_REGISTER = 8'h00;
parameter [7:0] PF0_CAPABILITY_POINTER = 8'h50;
parameter [23:0] PF0_CLASS_CODE = 24'h000000;
parameter [15:0] PF0_DEVICE_ID = 16'h0000;
parameter PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT = "TRUE";
parameter PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
parameter PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
parameter PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE = "TRUE";
parameter PF0_DEV_CAP2_LTR_SUPPORT = "TRUE";
parameter [1:0] PF0_DEV_CAP2_OBFF_SUPPORT = 2'h0;
parameter PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT = "FALSE";
parameter PF0_DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
parameter PF0_DEV_CAP_ENDPOINT_L1_LATENCY = 0;
parameter PF0_DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
parameter PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "TRUE";
parameter [2:0] PF0_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
parameter [11:0] PF0_DPA_CAP_NEXTPTR = 12'h000;
parameter [4:0] PF0_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
parameter PF0_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
parameter [3:0] PF0_DPA_CAP_VER = 4'h1;
parameter [11:0] PF0_DSN_CAP_NEXTPTR = 12'h10C;
parameter [4:0] PF0_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
parameter PF0_EXPANSION_ROM_ENABLE = "FALSE";
parameter [7:0] PF0_INTERRUPT_LINE = 8'h00;
parameter [2:0] PF0_INTERRUPT_PIN = 3'h1;
parameter PF0_LINK_CAP_ASPM_SUPPORT = 0;
parameter PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
parameter PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
parameter PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 = 7;
parameter PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
parameter PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
parameter PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 = 7;
parameter PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
parameter PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
parameter PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 = 7;
parameter PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
parameter PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
parameter PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 = 7;
parameter PF0_LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
parameter [9:0] PF0_LTR_CAP_MAX_NOSNOOP_LAT = 10'h000;
parameter [9:0] PF0_LTR_CAP_MAX_SNOOP_LAT = 10'h000;
parameter [11:0] PF0_LTR_CAP_NEXTPTR = 12'h000;
parameter [3:0] PF0_LTR_CAP_VER = 4'h1;
parameter [7:0] PF0_MSIX_CAP_NEXTPTR = 8'h00;
parameter PF0_MSIX_CAP_PBA_BIR = 0;
parameter [28:0] PF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
parameter PF0_MSIX_CAP_TABLE_BIR = 0;
parameter [28:0] PF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
parameter [10:0] PF0_MSIX_CAP_TABLE_SIZE = 11'h000;
parameter PF0_MSI_CAP_MULTIMSGCAP = 0;
parameter [7:0] PF0_MSI_CAP_NEXTPTR = 8'h00;
parameter [11:0] PF0_PB_CAP_NEXTPTR = 12'h000;
parameter PF0_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
parameter [3:0] PF0_PB_CAP_VER = 4'h1;
parameter [7:0] PF0_PM_CAP_ID = 8'h01;
parameter [7:0] PF0_PM_CAP_NEXTPTR = 8'h00;
parameter PF0_PM_CAP_PMESUPPORT_D0 = "TRUE";
parameter PF0_PM_CAP_PMESUPPORT_D1 = "TRUE";
parameter PF0_PM_CAP_PMESUPPORT_D3HOT = "TRUE";
parameter PF0_PM_CAP_SUPP_D1_STATE = "TRUE";
parameter [2:0] PF0_PM_CAP_VER_ID = 3'h3;
parameter PF0_PM_CSR_NOSOFTRESET = "TRUE";
parameter PF0_RBAR_CAP_ENABLE = "FALSE";
parameter [2:0] PF0_RBAR_CAP_INDEX0 = 3'h0;
parameter [2:0] PF0_RBAR_CAP_INDEX1 = 3'h0;
parameter [2:0] PF0_RBAR_CAP_INDEX2 = 3'h0;
parameter [11:0] PF0_RBAR_CAP_NEXTPTR = 12'h000;
parameter [19:0] PF0_RBAR_CAP_SIZE0 = 20'h00000;
parameter [19:0] PF0_RBAR_CAP_SIZE1 = 20'h00000;
parameter [19:0] PF0_RBAR_CAP_SIZE2 = 20'h00000;
parameter [3:0] PF0_RBAR_CAP_VER = 4'h1;
parameter [2:0] PF0_RBAR_NUM = 3'h1;
parameter [7:0] PF0_REVISION_ID = 8'h00;
parameter [4:0] PF0_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
parameter [2:0] PF0_SRIOV_BAR0_CONTROL = 3'h4;
parameter [4:0] PF0_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
parameter [2:0] PF0_SRIOV_BAR1_CONTROL = 3'h0;
parameter [4:0] PF0_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
parameter [2:0] PF0_SRIOV_BAR2_CONTROL = 3'h4;
parameter [4:0] PF0_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
parameter [2:0] PF0_SRIOV_BAR3_CONTROL = 3'h0;
parameter [4:0] PF0_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
parameter [2:0] PF0_SRIOV_BAR4_CONTROL = 3'h4;
parameter [4:0] PF0_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
parameter [2:0] PF0_SRIOV_BAR5_CONTROL = 3'h0;
parameter [15:0] PF0_SRIOV_CAP_INITIAL_VF = 16'h0000;
parameter [11:0] PF0_SRIOV_CAP_NEXTPTR = 12'h000;
parameter [15:0] PF0_SRIOV_CAP_TOTAL_VF = 16'h0000;
parameter [3:0] PF0_SRIOV_CAP_VER = 4'h1;
parameter [15:0] PF0_SRIOV_FIRST_VF_OFFSET = 16'h0000;
parameter [15:0] PF0_SRIOV_FUNC_DEP_LINK = 16'h0000;
parameter [31:0] PF0_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
parameter [15:0] PF0_SRIOV_VF_DEVICE_ID = 16'h0000;
parameter [15:0] PF0_SUBSYSTEM_ID = 16'h0000;
parameter PF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
parameter PF0_TPHR_CAP_ENABLE = "FALSE";
parameter PF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
parameter [11:0] PF0_TPHR_CAP_NEXTPTR = 12'h000;
parameter [2:0] PF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
parameter [1:0] PF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
parameter [10:0] PF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
parameter [3:0] PF0_TPHR_CAP_VER = 4'h1;
parameter [11:0] PF0_VC_CAP_NEXTPTR = 12'h000;
parameter [3:0] PF0_VC_CAP_VER = 4'h1;
parameter PF1_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
parameter PF1_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
parameter [11:0] PF1_AER_CAP_NEXTPTR = 12'h000;
parameter [11:0] PF1_ARI_CAP_NEXTPTR = 12'h000;
parameter [7:0] PF1_ARI_CAP_NEXT_FUNC = 8'h00;
parameter [4:0] PF1_BAR0_APERTURE_SIZE = 5'h03;
parameter [2:0] PF1_BAR0_CONTROL = 3'h4;
parameter [4:0] PF1_BAR1_APERTURE_SIZE = 5'h00;
parameter [2:0] PF1_BAR1_CONTROL = 3'h0;
parameter [4:0] PF1_BAR2_APERTURE_SIZE = 5'h03;
parameter [2:0] PF1_BAR2_CONTROL = 3'h4;
parameter [4:0] PF1_BAR3_APERTURE_SIZE = 5'h03;
parameter [2:0] PF1_BAR3_CONTROL = 3'h0;
parameter [4:0] PF1_BAR4_APERTURE_SIZE = 5'h03;
parameter [2:0] PF1_BAR4_CONTROL = 3'h4;
parameter [4:0] PF1_BAR5_APERTURE_SIZE = 5'h03;
parameter [2:0] PF1_BAR5_CONTROL = 3'h0;
parameter [7:0] PF1_BIST_REGISTER = 8'h00;
parameter [7:0] PF1_CAPABILITY_POINTER = 8'h50;
parameter [23:0] PF1_CLASS_CODE = 24'h000000;
parameter [15:0] PF1_DEVICE_ID = 16'h0000;
parameter [2:0] PF1_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
parameter [11:0] PF1_DPA_CAP_NEXTPTR = 12'h000;
parameter [4:0] PF1_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
parameter PF1_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
parameter [3:0] PF1_DPA_CAP_VER = 4'h1;
parameter [11:0] PF1_DSN_CAP_NEXTPTR = 12'h10C;
parameter [4:0] PF1_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
parameter PF1_EXPANSION_ROM_ENABLE = "FALSE";
parameter [7:0] PF1_INTERRUPT_LINE = 8'h00;
parameter [2:0] PF1_INTERRUPT_PIN = 3'h1;
parameter [7:0] PF1_MSIX_CAP_NEXTPTR = 8'h00;
parameter PF1_MSIX_CAP_PBA_BIR = 0;
parameter [28:0] PF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
parameter PF1_MSIX_CAP_TABLE_BIR = 0;
parameter [28:0] PF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
parameter [10:0] PF1_MSIX_CAP_TABLE_SIZE = 11'h000;
parameter PF1_MSI_CAP_MULTIMSGCAP = 0;
parameter [7:0] PF1_MSI_CAP_NEXTPTR = 8'h00;
parameter [11:0] PF1_PB_CAP_NEXTPTR = 12'h000;
parameter PF1_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
parameter [3:0] PF1_PB_CAP_VER = 4'h1;
parameter [7:0] PF1_PM_CAP_ID = 8'h01;
parameter [7:0] PF1_PM_CAP_NEXTPTR = 8'h00;
parameter [2:0] PF1_PM_CAP_VER_ID = 3'h3;
parameter PF1_RBAR_CAP_ENABLE = "FALSE";
parameter [2:0] PF1_RBAR_CAP_INDEX0 = 3'h0;
parameter [2:0] PF1_RBAR_CAP_INDEX1 = 3'h0;
parameter [2:0] PF1_RBAR_CAP_INDEX2 = 3'h0;
parameter [11:0] PF1_RBAR_CAP_NEXTPTR = 12'h000;
parameter [19:0] PF1_RBAR_CAP_SIZE0 = 20'h00000;
parameter [19:0] PF1_RBAR_CAP_SIZE1 = 20'h00000;
parameter [19:0] PF1_RBAR_CAP_SIZE2 = 20'h00000;
parameter [3:0] PF1_RBAR_CAP_VER = 4'h1;
parameter [2:0] PF1_RBAR_NUM = 3'h1;
parameter [7:0] PF1_REVISION_ID = 8'h00;
parameter [4:0] PF1_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
parameter [2:0] PF1_SRIOV_BAR0_CONTROL = 3'h4;
parameter [4:0] PF1_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
parameter [2:0] PF1_SRIOV_BAR1_CONTROL = 3'h0;
parameter [4:0] PF1_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
parameter [2:0] PF1_SRIOV_BAR2_CONTROL = 3'h4;
parameter [4:0] PF1_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
parameter [2:0] PF1_SRIOV_BAR3_CONTROL = 3'h0;
parameter [4:0] PF1_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
parameter [2:0] PF1_SRIOV_BAR4_CONTROL = 3'h4;
parameter [4:0] PF1_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
parameter [2:0] PF1_SRIOV_BAR5_CONTROL = 3'h0;
parameter [15:0] PF1_SRIOV_CAP_INITIAL_VF = 16'h0000;
parameter [11:0] PF1_SRIOV_CAP_NEXTPTR = 12'h000;
parameter [15:0] PF1_SRIOV_CAP_TOTAL_VF = 16'h0000;
parameter [3:0] PF1_SRIOV_CAP_VER = 4'h1;
parameter [15:0] PF1_SRIOV_FIRST_VF_OFFSET = 16'h0000;
parameter [15:0] PF1_SRIOV_FUNC_DEP_LINK = 16'h0000;
parameter [31:0] PF1_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
parameter [15:0] PF1_SRIOV_VF_DEVICE_ID = 16'h0000;
parameter [15:0] PF1_SUBSYSTEM_ID = 16'h0000;
parameter PF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
parameter PF1_TPHR_CAP_ENABLE = "FALSE";
parameter PF1_TPHR_CAP_INT_VEC_MODE = "TRUE";
parameter [11:0] PF1_TPHR_CAP_NEXTPTR = 12'h000;
parameter [2:0] PF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
parameter [1:0] PF1_TPHR_CAP_ST_TABLE_LOC = 2'h0;
parameter [10:0] PF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
parameter [3:0] PF1_TPHR_CAP_VER = 4'h1;
parameter PL_DISABLE_EI_INFER_IN_L0 = "FALSE";
parameter PL_DISABLE_GEN3_DC_BALANCE = "FALSE";
parameter PL_DISABLE_SCRAMBLING = "FALSE";
parameter PL_DISABLE_UPCONFIG_CAPABLE = "FALSE";
parameter PL_EQ_ADAPT_DISABLE_COEFF_CHECK = "FALSE";
parameter PL_EQ_ADAPT_DISABLE_PRESET_CHECK = "FALSE";
parameter [4:0] PL_EQ_ADAPT_ITER_COUNT = 5'h02;
parameter [1:0] PL_EQ_ADAPT_REJECT_RETRY_COUNT = 2'h1;
parameter PL_EQ_BYPASS_PHASE23 = "FALSE";
parameter PL_EQ_SHORT_ADAPT_PHASE = "FALSE";
parameter [15:0] PL_LANE0_EQ_CONTROL = 16'h3F00;
parameter [15:0] PL_LANE1_EQ_CONTROL = 16'h3F00;
parameter [15:0] PL_LANE2_EQ_CONTROL = 16'h3F00;
parameter [15:0] PL_LANE3_EQ_CONTROL = 16'h3F00;
parameter [15:0] PL_LANE4_EQ_CONTROL = 16'h3F00;
parameter [15:0] PL_LANE5_EQ_CONTROL = 16'h3F00;
parameter [15:0] PL_LANE6_EQ_CONTROL = 16'h3F00;
parameter [15:0] PL_LANE7_EQ_CONTROL = 16'h3F00;
parameter [2:0] PL_LINK_CAP_MAX_LINK_SPEED = 3'h4;
parameter [3:0] PL_LINK_CAP_MAX_LINK_WIDTH = 4'h8;
parameter PL_N_FTS_COMCLK_GEN1 = 255;
parameter PL_N_FTS_COMCLK_GEN2 = 255;
parameter PL_N_FTS_COMCLK_GEN3 = 255;
parameter PL_N_FTS_GEN1 = 255;
parameter PL_N_FTS_GEN2 = 255;
parameter PL_N_FTS_GEN3 = 255;
parameter PL_SIM_FAST_LINK_TRAINING = "FALSE";
parameter PL_UPSTREAM_FACING = "TRUE";
parameter [15:0] PM_ASPML0S_TIMEOUT = 16'h05DC;
parameter [19:0] PM_ASPML1_ENTRY_DELAY = 20'h00000;
parameter PM_ENABLE_SLOT_POWER_CAPTURE = "TRUE";
parameter [31:0] PM_L1_REENTRY_DELAY = 32'h00000000;
parameter [19:0] PM_PME_SERVICE_TIMEOUT_DELAY = 20'h186A0;
parameter [15:0] PM_PME_TURNOFF_ACK_DELAY = 16'h0064;
parameter SIM_VERSION = "1.0";
parameter SPARE_BIT0 = 0;
parameter SPARE_BIT1 = 0;
parameter SPARE_BIT2 = 0;
parameter SPARE_BIT3 = 0;
parameter SPARE_BIT4 = 0;
parameter SPARE_BIT5 = 0;
parameter SPARE_BIT6 = 0;
parameter SPARE_BIT7 = 0;
parameter SPARE_BIT8 = 0;
parameter [7:0] SPARE_BYTE0 = 8'h00;
parameter [7:0] SPARE_BYTE1 = 8'h00;
parameter [7:0] SPARE_BYTE2 = 8'h00;
parameter [7:0] SPARE_BYTE3 = 8'h00;
parameter [31:0] SPARE_WORD0 = 32'h00000000;
parameter [31:0] SPARE_WORD1 = 32'h00000000;
parameter [31:0] SPARE_WORD2 = 32'h00000000;
parameter [31:0] SPARE_WORD3 = 32'h00000000;
parameter SRIOV_CAP_ENABLE = "FALSE";
parameter [23:0] TL_COMPL_TIMEOUT_REG0 = 24'hBEBC20;
parameter [27:0] TL_COMPL_TIMEOUT_REG1 = 28'h0000000;
parameter [11:0] TL_CREDITS_CD = 12'h3E0;
parameter [7:0] TL_CREDITS_CH = 8'h20;
parameter [11:0] TL_CREDITS_NPD = 12'h028;
parameter [7:0] TL_CREDITS_NPH = 8'h20;
parameter [11:0] TL_CREDITS_PD = 12'h198;
parameter [7:0] TL_CREDITS_PH = 8'h20;
parameter TL_ENABLE_MESSAGE_RID_CHECK_ENABLE = "TRUE";
parameter TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
parameter TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
parameter TL_LEGACY_MODE_ENABLE = "FALSE";
parameter TL_PF_ENABLE_REG = "FALSE";
parameter TL_TAG_MGMT_ENABLE = "TRUE";
parameter [11:0] VF0_ARI_CAP_NEXTPTR = 12'h000;
parameter [7:0] VF0_CAPABILITY_POINTER = 8'h50;
parameter VF0_MSIX_CAP_PBA_BIR = 0;
parameter [28:0] VF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
parameter VF0_MSIX_CAP_TABLE_BIR = 0;
parameter [28:0] VF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
parameter [10:0] VF0_MSIX_CAP_TABLE_SIZE = 11'h000;
parameter VF0_MSI_CAP_MULTIMSGCAP = 0;
parameter [7:0] VF0_PM_CAP_ID = 8'h01;
parameter [7:0] VF0_PM_CAP_NEXTPTR = 8'h00;
parameter [2:0] VF0_PM_CAP_VER_ID = 3'h3;
parameter VF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
parameter VF0_TPHR_CAP_ENABLE = "FALSE";
parameter VF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
parameter [11:0] VF0_TPHR_CAP_NEXTPTR = 12'h000;
parameter [2:0] VF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
parameter [1:0] VF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
parameter [10:0] VF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
parameter [3:0] VF0_TPHR_CAP_VER = 4'h1;
parameter [11:0] VF1_ARI_CAP_NEXTPTR = 12'h000;
parameter VF1_MSIX_CAP_PBA_BIR = 0;
parameter [28:0] VF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
parameter VF1_MSIX_CAP_TABLE_BIR = 0;
parameter [28:0] VF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
parameter [10:0] VF1_MSIX_CAP_TABLE_SIZE = 11'h000;
parameter VF1_MSI_CAP_MULTIMSGCAP = 0;
parameter [7:0] VF1_PM_CAP_ID = 8'h01;
parameter [7:0] VF1_PM_CAP_NEXTPTR = 8'h00;
parameter [2:0] VF1_PM_CAP_VER_ID = 3'h3;
parameter VF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
parameter VF1_TPHR_CAP_ENABLE = "FALSE";
parameter VF1_TPHR_CAP_INT_VEC_MODE = "TRUE";
parameter [11:0] VF1_TPHR_CAP_NEXTPTR = 12'h000;
parameter [2:0] VF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
parameter [1:0] VF1_TPHR_CAP_ST_TABLE_LOC = 2'h0;
parameter [10:0] VF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
parameter [3:0] VF1_TPHR_CAP_VER = 4'h1;
parameter [11:0] VF2_ARI_CAP_NEXTPTR = 12'h000;
parameter VF2_MSIX_CAP_PBA_BIR = 0;
parameter [28:0] VF2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
parameter VF2_MSIX_CAP_TABLE_BIR = 0;
parameter [28:0] VF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
parameter [10:0] VF2_MSIX_CAP_TABLE_SIZE = 11'h000;
parameter VF2_MSI_CAP_MULTIMSGCAP = 0;
parameter [7:0] VF2_PM_CAP_ID = 8'h01;
parameter [7:0] VF2_PM_CAP_NEXTPTR = 8'h00;
parameter [2:0] VF2_PM_CAP_VER_ID = 3'h3;
parameter VF2_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
parameter VF2_TPHR_CAP_ENABLE = "FALSE";
parameter VF2_TPHR_CAP_INT_VEC_MODE = "TRUE";
parameter [11:0] VF2_TPHR_CAP_NEXTPTR = 12'h000;
parameter [2:0] VF2_TPHR_CAP_ST_MODE_SEL = 3'h0;
parameter [1:0] VF2_TPHR_CAP_ST_TABLE_LOC = 2'h0;
parameter [10:0] VF2_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
parameter [3:0] VF2_TPHR_CAP_VER = 4'h1;
parameter [11:0] VF3_ARI_CAP_NEXTPTR = 12'h000;
parameter VF3_MSIX_CAP_PBA_BIR = 0;
parameter [28:0] VF3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
parameter VF3_MSIX_CAP_TABLE_BIR = 0;
parameter [28:0] VF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
parameter [10:0] VF3_MSIX_CAP_TABLE_SIZE = 11'h000;
parameter VF3_MSI_CAP_MULTIMSGCAP = 0;
parameter [7:0] VF3_PM_CAP_ID = 8'h01;
parameter [7:0] VF3_PM_CAP_NEXTPTR = 8'h00;
parameter [2:0] VF3_PM_CAP_VER_ID = 3'h3;
parameter VF3_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
parameter VF3_TPHR_CAP_ENABLE = "FALSE";
parameter VF3_TPHR_CAP_INT_VEC_MODE = "TRUE";
parameter [11:0] VF3_TPHR_CAP_NEXTPTR = 12'h000;
parameter [2:0] VF3_TPHR_CAP_ST_MODE_SEL = 3'h0;
parameter [1:0] VF3_TPHR_CAP_ST_TABLE_LOC = 2'h0;
parameter [10:0] VF3_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
parameter [3:0] VF3_TPHR_CAP_VER = 4'h1;
parameter [11:0] VF4_ARI_CAP_NEXTPTR = 12'h000;
parameter VF4_MSIX_CAP_PBA_BIR = 0;
parameter [28:0] VF4_MSIX_CAP_PBA_OFFSET = 29'h00000050;
parameter VF4_MSIX_CAP_TABLE_BIR = 0;
parameter [28:0] VF4_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
parameter [10:0] VF4_MSIX_CAP_TABLE_SIZE = 11'h000;
parameter VF4_MSI_CAP_MULTIMSGCAP = 0;
parameter [7:0] VF4_PM_CAP_ID = 8'h01;
parameter [7:0] VF4_PM_CAP_NEXTPTR = 8'h00;
parameter [2:0] VF4_PM_CAP_VER_ID = 3'h3;
parameter VF4_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
parameter VF4_TPHR_CAP_ENABLE = "FALSE";
parameter VF4_TPHR_CAP_INT_VEC_MODE = "TRUE";
parameter [11:0] VF4_TPHR_CAP_NEXTPTR = 12'h000;
parameter [2:0] VF4_TPHR_CAP_ST_MODE_SEL = 3'h0;
parameter [1:0] VF4_TPHR_CAP_ST_TABLE_LOC = 2'h0;
parameter [10:0] VF4_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
parameter [3:0] VF4_TPHR_CAP_VER = 4'h1;
parameter [11:0] VF5_ARI_CAP_NEXTPTR = 12'h000;
parameter VF5_MSIX_CAP_PBA_BIR = 0;
parameter [28:0] VF5_MSIX_CAP_PBA_OFFSET = 29'h00000050;
parameter VF5_MSIX_CAP_TABLE_BIR = 0;
parameter [28:0] VF5_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
parameter [10:0] VF5_MSIX_CAP_TABLE_SIZE = 11'h000;
parameter VF5_MSI_CAP_MULTIMSGCAP = 0;
parameter [7:0] VF5_PM_CAP_ID = 8'h01;
parameter [7:0] VF5_PM_CAP_NEXTPTR = 8'h00;
parameter [2:0] VF5_PM_CAP_VER_ID = 3'h3;
parameter VF5_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
parameter VF5_TPHR_CAP_ENABLE = "FALSE";
parameter VF5_TPHR_CAP_INT_VEC_MODE = "TRUE";
parameter [11:0] VF5_TPHR_CAP_NEXTPTR = 12'h000;
parameter [2:0] VF5_TPHR_CAP_ST_MODE_SEL = 3'h0;
parameter [1:0] VF5_TPHR_CAP_ST_TABLE_LOC = 2'h0;
parameter [10:0] VF5_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
parameter [3:0] VF5_TPHR_CAP_VER = 4'h1;
endmodule
//#### END MODULE DEFINITION FOR: PCIE_3_0 ####

//#### BEGIN MODULE DEFINITION FOR :PCIE_A1 ###
module PCIE_A1 (
  CFGBUSNUMBER,
  CFGCOMMANDBUSMASTERENABLE,
  CFGCOMMANDINTERRUPTDISABLE,
  CFGCOMMANDIOENABLE,
  CFGCOMMANDMEMENABLE,
  CFGCOMMANDSERREN,
  CFGDEVCONTROLAUXPOWEREN,
  CFGDEVCONTROLCORRERRREPORTINGEN,
  CFGDEVCONTROLENABLERO,
  CFGDEVCONTROLEXTTAGEN,
  CFGDEVCONTROLFATALERRREPORTINGEN,
  CFGDEVCONTROLMAXPAYLOAD,
  CFGDEVCONTROLMAXREADREQ,
  CFGDEVCONTROLNONFATALREPORTINGEN,
  CFGDEVCONTROLNOSNOOPEN,
  CFGDEVCONTROLPHANTOMEN,
  CFGDEVCONTROLURERRREPORTINGEN,
  CFGDEVICENUMBER,
  CFGDEVSTATUSCORRERRDETECTED,
  CFGDEVSTATUSFATALERRDETECTED,
  CFGDEVSTATUSNONFATALERRDETECTED,
  CFGDEVSTATUSURDETECTED,
  CFGDO,
  CFGERRCPLRDYN,
  CFGFUNCTIONNUMBER,
  CFGINTERRUPTDO,
  CFGINTERRUPTMMENABLE,
  CFGINTERRUPTMSIENABLE,
  CFGINTERRUPTRDYN,
  CFGLINKCONTOLRCB,
  CFGLINKCONTROLASPMCONTROL,
  CFGLINKCONTROLCOMMONCLOCK,
  CFGLINKCONTROLEXTENDEDSYNC,
  CFGLTSSMSTATE,
  CFGPCIELINKSTATEN,
  CFGRDWRDONEN,
  CFGTOTURNOFFN,
  DBGBADDLLPSTATUS,
  DBGBADTLPLCRC,
  DBGBADTLPSEQNUM,
  DBGBADTLPSTATUS,
  DBGDLPROTOCOLSTATUS,
  DBGFCPROTOCOLERRSTATUS,
  DBGMLFRMDLENGTH,
  DBGMLFRMDMPS,
  DBGMLFRMDTCVC,
  DBGMLFRMDTLPSTATUS,
  DBGMLFRMDUNRECTYPE,
  DBGPOISTLPSTATUS,
  DBGRCVROVERFLOWSTATUS,
  DBGREGDETECTEDCORRECTABLE,
  DBGREGDETECTEDFATAL,
  DBGREGDETECTEDNONFATAL,
  DBGREGDETECTEDUNSUPPORTED,
  DBGRPLYROLLOVERSTATUS,
  DBGRPLYTIMEOUTSTATUS,
  DBGURNOBARHIT,
  DBGURPOISCFGWR,
  DBGURSTATUS,
  DBGURUNSUPMSG,
  MIMRXRADDR,
  MIMRXREN,
  MIMRXWADDR,
  MIMRXWDATA,
  MIMRXWEN,
  MIMTXRADDR,
  MIMTXREN,
  MIMTXWADDR,
  MIMTXWDATA,
  MIMTXWEN,
  PIPEGTPOWERDOWNA,
  PIPEGTPOWERDOWNB,
  PIPEGTTXELECIDLEA,
  PIPEGTTXELECIDLEB,
  PIPERXPOLARITYA,
  PIPERXPOLARITYB,
  PIPERXRESETA,
  PIPERXRESETB,
  PIPETXCHARDISPMODEA,
  PIPETXCHARDISPMODEB,
  PIPETXCHARDISPVALA,
  PIPETXCHARDISPVALB,
  PIPETXCHARISKA,
  PIPETXCHARISKB,
  PIPETXDATAA,
  PIPETXDATAB,
  PIPETXRCVRDETA,
  PIPETXRCVRDETB,
  RECEIVEDHOTRESET,
  TRNFCCPLD,
  TRNFCCPLH,
  TRNFCNPD,
  TRNFCNPH,
  TRNFCPD,
  TRNFCPH,
  TRNLNKUPN,
  TRNRBARHITN,
  TRNRD,
  TRNREOFN,
  TRNRERRFWDN,
  TRNRSOFN,
  TRNRSRCDSCN,
  TRNRSRCRDYN,
  TRNTBUFAV,
  TRNTCFGREQN,
  TRNTDSTRDYN,
  TRNTERRDROPN,
  USERRSTN,
  CFGDEVID,
  CFGDSN,
  CFGDWADDR,
  CFGERRCORN,
  CFGERRCPLABORTN,
  CFGERRCPLTIMEOUTN,
  CFGERRECRCN,
  CFGERRLOCKEDN,
  CFGERRPOSTEDN,
  CFGERRTLPCPLHEADER,
  CFGERRURN,
  CFGINTERRUPTASSERTN,
  CFGINTERRUPTDI,
  CFGINTERRUPTN,
  CFGPMWAKEN,
  CFGRDENN,
  CFGREVID,
  CFGSUBSYSID,
  CFGSUBSYSVENID,
  CFGTRNPENDINGN,
  CFGTURNOFFOKN,
  CFGVENID,
  CLOCKLOCKED,
  MGTCLK,
  MIMRXRDATA,
  MIMTXRDATA,
  PIPEGTRESETDONEA,
  PIPEGTRESETDONEB,
  PIPEPHYSTATUSA,
  PIPEPHYSTATUSB,
  PIPERXCHARISKA,
  PIPERXCHARISKB,
  PIPERXDATAA,
  PIPERXDATAB,
  PIPERXENTERELECIDLEA,
  PIPERXENTERELECIDLEB,
  PIPERXSTATUSA,
  PIPERXSTATUSB,
  SYSRESETN,
  TRNFCSEL,
  TRNRDSTRDYN,
  TRNRNPOKN,
  TRNTCFGGNTN,
  TRNTD,
  TRNTEOFN,
  TRNTERRFWDN,
  TRNTSOFN,
  TRNTSRCDSCN,
  TRNTSRCRDYN,
  TRNTSTRN,
  USERCLK
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CFGERRCORN ;
input CFGERRCPLABORTN ;
input CFGERRCPLTIMEOUTN ;
input CFGERRECRCN ;
input CFGERRLOCKEDN ;
input CFGERRPOSTEDN ;
input CFGERRURN ;
input CFGINTERRUPTASSERTN ;
input CFGINTERRUPTN ;
input CFGPMWAKEN ;
input CFGRDENN ;
input CFGTRNPENDINGN ;
input CFGTURNOFFOKN ;
input CLOCKLOCKED ;
input MGTCLK ;
input PIPEGTRESETDONEA ;
input PIPEGTRESETDONEB ;
input PIPEPHYSTATUSA ;
input PIPEPHYSTATUSB ;
input PIPERXENTERELECIDLEA ;
input PIPERXENTERELECIDLEB ;
input SYSRESETN ;
input TRNRDSTRDYN ;
input TRNRNPOKN ;
input TRNTCFGGNTN ;
input TRNTEOFN ;
input TRNTERRFWDN ;
input TRNTSOFN ;
input TRNTSRCDSCN ;
input TRNTSRCRDYN ;
input TRNTSTRN ;
input USERCLK ;
input [15:0] CFGDEVID ;
input [15:0] CFGSUBSYSID ;
input [15:0] CFGSUBSYSVENID ;
input [15:0] CFGVENID ;
input [15:0] PIPERXDATAA ;
input [15:0] PIPERXDATAB ;
input [1:0] PIPERXCHARISKA ;
input [1:0] PIPERXCHARISKB ;
input [2:0] PIPERXSTATUSA ;
input [2:0] PIPERXSTATUSB ;
input [2:0] TRNFCSEL ;
input [31:0] TRNTD ;
input [34:0] MIMRXRDATA ;
input [35:0] MIMTXRDATA ;
input [47:0] CFGERRTLPCPLHEADER ;
input [63:0] CFGDSN ;
input [7:0] CFGINTERRUPTDI ;
input [7:0] CFGREVID ;
input [9:0] CFGDWADDR ;
output CFGCOMMANDBUSMASTERENABLE ;
output CFGCOMMANDINTERRUPTDISABLE ;
output CFGCOMMANDIOENABLE ;
output CFGCOMMANDMEMENABLE ;
output CFGCOMMANDSERREN ;
output CFGDEVCONTROLAUXPOWEREN ;
output CFGDEVCONTROLCORRERRREPORTINGEN ;
output CFGDEVCONTROLENABLERO ;
output CFGDEVCONTROLEXTTAGEN ;
output CFGDEVCONTROLFATALERRREPORTINGEN ;
output CFGDEVCONTROLNONFATALREPORTINGEN ;
output CFGDEVCONTROLNOSNOOPEN ;
output CFGDEVCONTROLPHANTOMEN ;
output CFGDEVCONTROLURERRREPORTINGEN ;
output CFGDEVSTATUSCORRERRDETECTED ;
output CFGDEVSTATUSFATALERRDETECTED ;
output CFGDEVSTATUSNONFATALERRDETECTED ;
output CFGDEVSTATUSURDETECTED ;
output CFGERRCPLRDYN ;
output CFGINTERRUPTMSIENABLE ;
output CFGINTERRUPTRDYN ;
output CFGLINKCONTOLRCB ;
output CFGLINKCONTROLCOMMONCLOCK ;
output CFGLINKCONTROLEXTENDEDSYNC ;
output CFGRDWRDONEN ;
output CFGTOTURNOFFN ;
output DBGBADDLLPSTATUS ;
output DBGBADTLPLCRC ;
output DBGBADTLPSEQNUM ;
output DBGBADTLPSTATUS ;
output DBGDLPROTOCOLSTATUS ;
output DBGFCPROTOCOLERRSTATUS ;
output DBGMLFRMDLENGTH ;
output DBGMLFRMDMPS ;
output DBGMLFRMDTCVC ;
output DBGMLFRMDTLPSTATUS ;
output DBGMLFRMDUNRECTYPE ;
output DBGPOISTLPSTATUS ;
output DBGRCVROVERFLOWSTATUS ;
output DBGREGDETECTEDCORRECTABLE ;
output DBGREGDETECTEDFATAL ;
output DBGREGDETECTEDNONFATAL ;
output DBGREGDETECTEDUNSUPPORTED ;
output DBGRPLYROLLOVERSTATUS ;
output DBGRPLYTIMEOUTSTATUS ;
output DBGURNOBARHIT ;
output DBGURPOISCFGWR ;
output DBGURSTATUS ;
output DBGURUNSUPMSG ;
output MIMRXREN ;
output MIMRXWEN ;
output MIMTXREN ;
output MIMTXWEN ;
output PIPEGTTXELECIDLEA ;
output PIPEGTTXELECIDLEB ;
output PIPERXPOLARITYA ;
output PIPERXPOLARITYB ;
output PIPERXRESETA ;
output PIPERXRESETB ;
output PIPETXRCVRDETA ;
output PIPETXRCVRDETB ;
output RECEIVEDHOTRESET ;
output TRNLNKUPN ;
output TRNREOFN ;
output TRNRERRFWDN ;
output TRNRSOFN ;
output TRNRSRCDSCN ;
output TRNRSRCRDYN ;
output TRNTCFGREQN ;
output TRNTDSTRDYN ;
output TRNTERRDROPN ;
output USERRSTN ;
output [11:0] MIMRXRADDR ;
output [11:0] MIMRXWADDR ;
output [11:0] MIMTXRADDR ;
output [11:0] MIMTXWADDR ;
output [11:0] TRNFCCPLD ;
output [11:0] TRNFCNPD ;
output [11:0] TRNFCPD ;
output [15:0] PIPETXDATAA ;
output [15:0] PIPETXDATAB ;
output [1:0] CFGLINKCONTROLASPMCONTROL ;
output [1:0] PIPEGTPOWERDOWNA ;
output [1:0] PIPEGTPOWERDOWNB ;
output [1:0] PIPETXCHARDISPMODEA ;
output [1:0] PIPETXCHARDISPMODEB ;
output [1:0] PIPETXCHARDISPVALA ;
output [1:0] PIPETXCHARDISPVALB ;
output [1:0] PIPETXCHARISKA ;
output [1:0] PIPETXCHARISKB ;
output [2:0] CFGDEVCONTROLMAXPAYLOAD ;
output [2:0] CFGDEVCONTROLMAXREADREQ ;
output [2:0] CFGFUNCTIONNUMBER ;
output [2:0] CFGINTERRUPTMMENABLE ;
output [2:0] CFGPCIELINKSTATEN ;
output [31:0] CFGDO ;
output [31:0] TRNRD ;
output [34:0] MIMRXWDATA ;
output [35:0] MIMTXWDATA ;
output [4:0] CFGDEVICENUMBER ;
output [4:0] CFGLTSSMSTATE ;
output [5:0] TRNTBUFAV ;
output [6:0] TRNRBARHITN ;
output [7:0] CFGBUSNUMBER ;
output [7:0] CFGINTERRUPTDO ;
output [7:0] TRNFCCPLH ;
output [7:0] TRNFCNPH ;
output [7:0] TRNFCPH ;
parameter [31:0] BAR0 = 32'h00000000;
parameter [31:0] BAR1 = 32'h00000000;
parameter [31:0] BAR2 = 32'h00000000;
parameter [31:0] BAR3 = 32'h00000000;
parameter [31:0] BAR4 = 32'h00000000;
parameter [31:0] BAR5 = 32'h00000000;
parameter [31:0] CARDBUS_CIS_POINTER = 32'h00000000;
parameter [23:0] CLASS_CODE = 24'h000000;
parameter DEV_CAP_ENDPOINT_L0S_LATENCY = 7;
parameter DEV_CAP_ENDPOINT_L1_LATENCY = 7;
parameter DEV_CAP_EXT_TAG_SUPPORTED = "FALSE";
parameter DEV_CAP_MAX_PAYLOAD_SUPPORTED = 2;
parameter DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT = 0;
parameter DEV_CAP_ROLE_BASED_ERROR = "TRUE";
parameter DISABLE_BAR_FILTERING = "FALSE";
parameter DISABLE_ID_CHECK = "FALSE";
parameter DISABLE_SCRAMBLING = "FALSE";
parameter ENABLE_RX_TD_ECRC_TRIM = "FALSE";
parameter [21:0] EXPANSION_ROM = 22'h000000;
parameter FAST_TRAIN = "FALSE";
parameter GTP_SEL = 0;
parameter LINK_CAP_ASPM_SUPPORT = 1;
parameter LINK_CAP_L0S_EXIT_LATENCY = 7;
parameter LINK_CAP_L1_EXIT_LATENCY = 7;
parameter LINK_STATUS_SLOT_CLOCK_CONFIG = "FALSE";
parameter [14:0] LL_ACK_TIMEOUT = 15'h0204;
parameter LL_ACK_TIMEOUT_EN = "FALSE";
parameter [14:0] LL_REPLAY_TIMEOUT = 15'h060D;
parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
parameter MSI_CAP_MULTIMSGCAP = 0;
parameter MSI_CAP_MULTIMSG_EXTENSION = 0;
parameter [3:0] PCIE_CAP_CAPABILITY_VERSION = 4'h1;
parameter [3:0] PCIE_CAP_DEVICE_PORT_TYPE = 4'h0;
parameter [4:0] PCIE_CAP_INT_MSG_NUM = 5'b00000;
parameter PCIE_CAP_SLOT_IMPLEMENTED = "FALSE";
parameter [11:0] PCIE_GENERIC = 12'h000;
parameter PLM_AUTO_CONFIG = "FALSE";
parameter PM_CAP_AUXCURRENT = 0;
parameter PM_CAP_D1SUPPORT = "TRUE";
parameter PM_CAP_D2SUPPORT = "TRUE";
parameter PM_CAP_DSI = "FALSE";
parameter [4:0] PM_CAP_PMESUPPORT = 5'b01111;
parameter PM_CAP_PME_CLOCK = "FALSE";
parameter PM_CAP_VERSION = 3;
parameter [7:0] PM_DATA0 = 8'h1E;
parameter [7:0] PM_DATA1 = 8'h1E;
parameter [7:0] PM_DATA2 = 8'h1E;
parameter [7:0] PM_DATA3 = 8'h1E;
parameter [7:0] PM_DATA4 = 8'h1E;
parameter [7:0] PM_DATA5 = 8'h1E;
parameter [7:0] PM_DATA6 = 8'h1E;
parameter [7:0] PM_DATA7 = 8'h1E;
parameter [1:0] PM_DATA_SCALE0 = 2'b01;
parameter [1:0] PM_DATA_SCALE1 = 2'b01;
parameter [1:0] PM_DATA_SCALE2 = 2'b01;
parameter [1:0] PM_DATA_SCALE3 = 2'b01;
parameter [1:0] PM_DATA_SCALE4 = 2'b01;
parameter [1:0] PM_DATA_SCALE5 = 2'b01;
parameter [1:0] PM_DATA_SCALE6 = 2'b01;
parameter [1:0] PM_DATA_SCALE7 = 2'b01;
parameter SIM_VERSION = "1.0";
parameter SLOT_CAP_ATT_BUTTON_PRESENT = "FALSE";
parameter SLOT_CAP_ATT_INDICATOR_PRESENT = "FALSE";
parameter SLOT_CAP_POWER_INDICATOR_PRESENT = "FALSE";
parameter TL_RX_RAM_RADDR_LATENCY = 1;
parameter TL_RX_RAM_RDATA_LATENCY = 2;
parameter TL_RX_RAM_WRITE_LATENCY = 0;
parameter TL_TFC_DISABLE = "FALSE";
parameter TL_TX_CHECKS_DISABLE = "FALSE";
parameter TL_TX_RAM_RADDR_LATENCY = 0;
parameter TL_TX_RAM_RDATA_LATENCY = 2;
parameter USR_CFG = "FALSE";
parameter USR_EXT_CFG = "FALSE";
parameter VC0_CPL_INFINITE = "TRUE";
parameter [11:0] VC0_RX_RAM_LIMIT = 12'h01E;
parameter VC0_TOTAL_CREDITS_CD = 104;
parameter VC0_TOTAL_CREDITS_CH = 36;
parameter VC0_TOTAL_CREDITS_NPH = 8;
parameter VC0_TOTAL_CREDITS_PD = 288;
parameter VC0_TOTAL_CREDITS_PH = 32;
parameter VC0_TX_LASTPACKET = 31;
endmodule
//#### END MODULE DEFINITION FOR: PCIE_A1 ####

//#### BEGIN MODULE DEFINITION FOR :PCIE_EP ###
module PCIE_EP (
	BUSMASTERENABLE,
	CRMDOHOTRESETN,
	CRMPWRSOFTRESETN,
	DLLTXPMDLLPOUTSTANDING,
	INTERRUPTDISABLE,
	IOSPACEENABLE,
	L0CFGLOOPBACKACK,
	L0COMPLETERID,
	L0DLLERRORVECTOR,
	L0DLLRXACKOUTSTANDING,
	L0DLLTXNONFCOUTSTANDING,
	L0DLLTXOUTSTANDING,
	L0DLLVCSTATUS,
	L0DLUPDOWN,
	L0FIRSTCFGWRITEOCCURRED,
	L0LTSSMSTATE,
	L0MACENTEREDL0,
	L0MACLINKTRAINING,
	L0MACLINKUP,
	L0MACNEGOTIATEDLINKWIDTH,
	L0MACNEWSTATEACK,
	L0MACRXL0SSTATE,
	L0MSIENABLE0,
	L0MULTIMSGEN0,
	L0PMEACK,
	L0PMEEN,
	L0PMEREQOUT,
	L0PWRL1STATE,
	L0PWRL23READYSTATE,
	L0PWRSTATE0,
	L0PWRTURNOFFREQ,
	L0PWRTXL0SSTATE,
	L0RXDLLPM,
	L0RXDLLPMTYPE,
	L0RXMACLINKERROR,
	L0STATSCFGOTHERRECEIVED,
	L0STATSCFGOTHERTRANSMITTED,
	L0STATSCFGRECEIVED,
	L0STATSCFGTRANSMITTED,
	L0STATSDLLPRECEIVED,
	L0STATSDLLPTRANSMITTED,
	L0STATSOSRECEIVED,
	L0STATSOSTRANSMITTED,
	L0STATSTLPRECEIVED,
	L0STATSTLPTRANSMITTED,
	L0UNLOCKRECEIVED,
	LLKRXCHCOMPLETIONAVAILABLEN,
	LLKRXCHNONPOSTEDAVAILABLEN,
	LLKRXCHPOSTEDAVAILABLEN,
	LLKRXDATA,
	LLKRXEOFN,
	LLKRXEOPN,
	LLKRXPREFERREDTYPE,
	LLKRXSOFN,
	LLKRXSOPN,
	LLKRXSRCLASTREQN,
	LLKRXSRCRDYN,
	LLKRXVALIDN,
	LLKTCSTATUS,
	LLKTXCHANSPACE,
	LLKTXCHCOMPLETIONREADYN,
	LLKTXCHNONPOSTEDREADYN,
	LLKTXCHPOSTEDREADYN,
	LLKTXCONFIGREADYN,
	LLKTXDSTRDYN,
	MAXPAYLOADSIZE,
	MAXREADREQUESTSIZE,
	MEMSPACEENABLE,
	MGMTPSO,
	MGMTRDATA,
	MGMTSTATSCREDIT,
	MIMDLLBRADD,
	MIMDLLBREN,
	MIMDLLBWADD,
	MIMDLLBWDATA,
	MIMDLLBWEN,
	MIMRXBRADD,
	MIMRXBREN,
	MIMRXBWADD,
	MIMRXBWDATA,
	MIMRXBWEN,
	MIMTXBRADD,
	MIMTXBREN,
	MIMTXBWADD,
	MIMTXBWDATA,
	MIMTXBWEN,
	PARITYERRORRESPONSE,
	PIPEDESKEWLANESL0,
	PIPEDESKEWLANESL1,
	PIPEDESKEWLANESL2,
	PIPEDESKEWLANESL3,
	PIPEDESKEWLANESL4,
	PIPEDESKEWLANESL5,
	PIPEDESKEWLANESL6,
	PIPEDESKEWLANESL7,
	PIPEPOWERDOWNL0,
	PIPEPOWERDOWNL1,
	PIPEPOWERDOWNL2,
	PIPEPOWERDOWNL3,
	PIPEPOWERDOWNL4,
	PIPEPOWERDOWNL5,
	PIPEPOWERDOWNL6,
	PIPEPOWERDOWNL7,
	PIPERESETL0,
	PIPERESETL1,
	PIPERESETL2,
	PIPERESETL3,
	PIPERESETL4,
	PIPERESETL5,
	PIPERESETL6,
	PIPERESETL7,
	PIPERXPOLARITYL0,
	PIPERXPOLARITYL1,
	PIPERXPOLARITYL2,
	PIPERXPOLARITYL3,
	PIPERXPOLARITYL4,
	PIPERXPOLARITYL5,
	PIPERXPOLARITYL6,
	PIPERXPOLARITYL7,
	PIPETXCOMPLIANCEL0,
	PIPETXCOMPLIANCEL1,
	PIPETXCOMPLIANCEL2,
	PIPETXCOMPLIANCEL3,
	PIPETXCOMPLIANCEL4,
	PIPETXCOMPLIANCEL5,
	PIPETXCOMPLIANCEL6,
	PIPETXCOMPLIANCEL7,
	PIPETXDATAKL0,
	PIPETXDATAKL1,
	PIPETXDATAKL2,
	PIPETXDATAKL3,
	PIPETXDATAKL4,
	PIPETXDATAKL5,
	PIPETXDATAKL6,
	PIPETXDATAKL7,
	PIPETXDATAL0,
	PIPETXDATAL1,
	PIPETXDATAL2,
	PIPETXDATAL3,
	PIPETXDATAL4,
	PIPETXDATAL5,
	PIPETXDATAL6,
	PIPETXDATAL7,
	PIPETXDETECTRXLOOPBACKL0,
	PIPETXDETECTRXLOOPBACKL1,
	PIPETXDETECTRXLOOPBACKL2,
	PIPETXDETECTRXLOOPBACKL3,
	PIPETXDETECTRXLOOPBACKL4,
	PIPETXDETECTRXLOOPBACKL5,
	PIPETXDETECTRXLOOPBACKL6,
	PIPETXDETECTRXLOOPBACKL7,
	PIPETXELECIDLEL0,
	PIPETXELECIDLEL1,
	PIPETXELECIDLEL2,
	PIPETXELECIDLEL3,
	PIPETXELECIDLEL4,
	PIPETXELECIDLEL5,
	PIPETXELECIDLEL6,
	PIPETXELECIDLEL7,
	SERRENABLE,
	URREPORTINGENABLE,

	AUXPOWER,
	COMPLIANCEAVOID,
	CRMCORECLK,
	CRMCORECLKDLO,
	CRMCORECLKRXO,
	CRMCORECLKTXO,
	CRMLINKRSTN,
	CRMMACRSTN,
	CRMMGMTRSTN,
	CRMNVRSTN,
	CRMURSTN,
	CRMUSERCFGRSTN,
	CRMUSERCLK,
	CRMUSERCLKRXO,
	CRMUSERCLKTXO,
	L0CFGDISABLESCRAMBLE,
	L0CFGLOOPBACKMASTER,
	L0LEGACYINTFUNCT0,
	L0MSIREQUEST0,
	L0PACKETHEADERFROMUSER,
	L0PMEREQIN,
	L0SETCOMPLETERABORTERROR,
	L0SETCOMPLETIONTIMEOUTCORRERROR,
	L0SETCOMPLETIONTIMEOUTUNCORRERROR,
	L0SETDETECTEDCORRERROR,
	L0SETDETECTEDFATALERROR,
	L0SETDETECTEDNONFATALERROR,
	L0SETUNEXPECTEDCOMPLETIONCORRERROR,
	L0SETUNEXPECTEDCOMPLETIONUNCORRERROR,
	L0SETUNSUPPORTEDREQUESTNONPOSTEDERROR,
	L0SETUNSUPPORTEDREQUESTOTHERERROR,
	L0SETUSERDETECTEDPARITYERROR,
	L0SETUSERMASTERDATAPARITY,
	L0SETUSERRECEIVEDMASTERABORT,
	L0SETUSERRECEIVEDTARGETABORT,
	L0SETUSERSIGNALLEDTARGETABORT,
	L0SETUSERSYSTEMERROR,
	L0TRANSACTIONSPENDING,
	LLKRXCHFIFO,
	LLKRXCHTC,
	LLKRXDSTCONTREQN,	
	LLKRXDSTREQN,
	LLKTXCHFIFO,
	LLKTXCHTC,
	LLKTXDATA,
	LLKTXENABLEN,
	LLKTXEOFN,
	LLKTXEOPN,
	LLKTXSOFN,
	LLKTXSOPN,
	LLKTXSRCDSCN,
	LLKTXSRCRDYN,
	MGMTADDR,
	MGMTBWREN,
	MGMTRDEN,
	MGMTSTATSCREDITSEL,
	MGMTWDATA,
	MGMTWREN,
	MIMDLLBRDATA,
	MIMRXBRDATA,
	MIMTXBRDATA,
	PIPEPHYSTATUSL0,
	PIPEPHYSTATUSL1,
	PIPEPHYSTATUSL2,
	PIPEPHYSTATUSL3,
	PIPEPHYSTATUSL4,
	PIPEPHYSTATUSL5,
	PIPEPHYSTATUSL6,
	PIPEPHYSTATUSL7,
	PIPERXCHANISALIGNEDL0,
	PIPERXCHANISALIGNEDL1,
	PIPERXCHANISALIGNEDL2,
	PIPERXCHANISALIGNEDL3,
	PIPERXCHANISALIGNEDL4,
	PIPERXCHANISALIGNEDL5,
	PIPERXCHANISALIGNEDL6,
	PIPERXCHANISALIGNEDL7,
	PIPERXDATAKL0,
	PIPERXDATAKL1,
	PIPERXDATAKL2,
	PIPERXDATAKL3,
	PIPERXDATAKL4,
	PIPERXDATAKL5,
	PIPERXDATAKL6,
	PIPERXDATAKL7,
	PIPERXDATAL0,
	PIPERXDATAL1,
	PIPERXDATAL2,
	PIPERXDATAL3,
	PIPERXDATAL4,
	PIPERXDATAL5,
	PIPERXDATAL6,
	PIPERXDATAL7,
	PIPERXELECIDLEL0,
	PIPERXELECIDLEL1,
	PIPERXELECIDLEL2,
	PIPERXELECIDLEL3,
	PIPERXELECIDLEL4,
	PIPERXELECIDLEL5,
	PIPERXELECIDLEL6,
	PIPERXELECIDLEL7,
	PIPERXSTATUSL0,
	PIPERXSTATUSL1,
	PIPERXSTATUSL2,
	PIPERXSTATUSL3,
	PIPERXSTATUSL4,
	PIPERXSTATUSL5,
	PIPERXSTATUSL6,
	PIPERXSTATUSL7,
	PIPERXVALIDL0,
	PIPERXVALIDL1,
	PIPERXVALIDL2,
	PIPERXVALIDL3,
	PIPERXVALIDL4,
	PIPERXVALIDL5,
	PIPERXVALIDL6,
	PIPERXVALIDL7

) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input AUXPOWER ;
input COMPLIANCEAVOID ;
input CRMCORECLK ;
input CRMCORECLKDLO ;
input CRMCORECLKRXO ;
input CRMCORECLKTXO ;
input CRMLINKRSTN ;
input CRMMACRSTN ;
input CRMMGMTRSTN ;
input CRMNVRSTN ;
input CRMURSTN ;
input CRMUSERCFGRSTN ;
input CRMUSERCLK ;
input CRMUSERCLKRXO ;
input CRMUSERCLKTXO ;
input L0CFGDISABLESCRAMBLE ;
input L0CFGLOOPBACKMASTER ;
input L0LEGACYINTFUNCT0 ;
input L0PMEREQIN ;
input L0SETCOMPLETERABORTERROR ;
input L0SETCOMPLETIONTIMEOUTCORRERROR ;
input L0SETCOMPLETIONTIMEOUTUNCORRERROR ;
input L0SETDETECTEDCORRERROR ;
input L0SETDETECTEDFATALERROR ;
input L0SETDETECTEDNONFATALERROR ;
input L0SETUNEXPECTEDCOMPLETIONCORRERROR ;
input L0SETUNEXPECTEDCOMPLETIONUNCORRERROR ;
input L0SETUNSUPPORTEDREQUESTNONPOSTEDERROR ;
input L0SETUNSUPPORTEDREQUESTOTHERERROR ;
input L0SETUSERDETECTEDPARITYERROR ;
input L0SETUSERMASTERDATAPARITY ;
input L0SETUSERRECEIVEDMASTERABORT ;
input L0SETUSERRECEIVEDTARGETABORT ;
input L0SETUSERSIGNALLEDTARGETABORT ;
input L0SETUSERSYSTEMERROR ;
input L0TRANSACTIONSPENDING ;
input LLKRXDSTCONTREQN ;
input LLKRXDSTREQN ;
input LLKTXEOFN ;
input LLKTXEOPN ;
input LLKTXSOFN ;
input LLKTXSOPN ;
input LLKTXSRCDSCN ;
input LLKTXSRCRDYN ;
input MGMTRDEN ;
input MGMTWREN ;
input PIPEPHYSTATUSL0 ;
input PIPEPHYSTATUSL1 ;
input PIPEPHYSTATUSL2 ;
input PIPEPHYSTATUSL3 ;
input PIPEPHYSTATUSL4 ;
input PIPEPHYSTATUSL5 ;
input PIPEPHYSTATUSL6 ;
input PIPEPHYSTATUSL7 ;
input PIPERXCHANISALIGNEDL0 ;
input PIPERXCHANISALIGNEDL1 ;
input PIPERXCHANISALIGNEDL2 ;
input PIPERXCHANISALIGNEDL3 ;
input PIPERXCHANISALIGNEDL4 ;
input PIPERXCHANISALIGNEDL5 ;
input PIPERXCHANISALIGNEDL6 ;
input PIPERXCHANISALIGNEDL7 ;
input PIPERXDATAKL0 ;
input PIPERXDATAKL1 ;
input PIPERXDATAKL2 ;
input PIPERXDATAKL3 ;
input PIPERXDATAKL4 ;
input PIPERXDATAKL5 ;
input PIPERXDATAKL6 ;
input PIPERXDATAKL7 ;
input PIPERXELECIDLEL0 ;
input PIPERXELECIDLEL1 ;
input PIPERXELECIDLEL2 ;
input PIPERXELECIDLEL3 ;
input PIPERXELECIDLEL4 ;
input PIPERXELECIDLEL5 ;
input PIPERXELECIDLEL6 ;
input PIPERXELECIDLEL7 ;
input PIPERXVALIDL0 ;
input PIPERXVALIDL1 ;
input PIPERXVALIDL2 ;
input PIPERXVALIDL3 ;
input PIPERXVALIDL4 ;
input PIPERXVALIDL5 ;
input PIPERXVALIDL6 ;
input PIPERXVALIDL7 ;
input [10:0] MGMTADDR ;
input [127:0] L0PACKETHEADERFROMUSER ;
input [1:0] LLKRXCHFIFO ;
input [1:0] LLKTXCHFIFO ;
input [1:0] LLKTXENABLEN ;
input [2:0] LLKRXCHTC ;
input [2:0] LLKTXCHTC ;
input [2:0] PIPERXSTATUSL0 ;
input [2:0] PIPERXSTATUSL1 ;
input [2:0] PIPERXSTATUSL2 ;
input [2:0] PIPERXSTATUSL3 ;
input [2:0] PIPERXSTATUSL4 ;
input [2:0] PIPERXSTATUSL5 ;
input [2:0] PIPERXSTATUSL6 ;
input [2:0] PIPERXSTATUSL7 ;
input [31:0] MGMTWDATA ;
input [3:0] L0MSIREQUEST0 ;
input [3:0] MGMTBWREN ;
input [63:0] LLKTXDATA ;
input [63:0] MIMDLLBRDATA ;
input [63:0] MIMRXBRDATA ;
input [63:0] MIMTXBRDATA ;
input [6:0] MGMTSTATSCREDITSEL ;
input [7:0] PIPERXDATAL0 ;
input [7:0] PIPERXDATAL1 ;
input [7:0] PIPERXDATAL2 ;
input [7:0] PIPERXDATAL3 ;
input [7:0] PIPERXDATAL4 ;
input [7:0] PIPERXDATAL5 ;
input [7:0] PIPERXDATAL6 ;
input [7:0] PIPERXDATAL7 ;
output BUSMASTERENABLE ;
output CRMDOHOTRESETN ;
output CRMPWRSOFTRESETN ;
output DLLTXPMDLLPOUTSTANDING ;
output INTERRUPTDISABLE ;
output IOSPACEENABLE ;
output L0CFGLOOPBACKACK ;
output L0DLLRXACKOUTSTANDING ;
output L0DLLTXNONFCOUTSTANDING ;
output L0DLLTXOUTSTANDING ;
output L0FIRSTCFGWRITEOCCURRED ;
output L0MACENTEREDL0 ;
output L0MACLINKTRAINING ;
output L0MACLINKUP ;
output L0MACNEWSTATEACK ;
output L0MACRXL0SSTATE ;
output L0MSIENABLE0 ;
output L0PMEACK ;
output L0PMEEN ;
output L0PMEREQOUT ;
output L0PWRL1STATE ;
output L0PWRL23READYSTATE ;
output L0PWRTURNOFFREQ ;
output L0PWRTXL0SSTATE ;
output L0RXDLLPM ;
output L0STATSCFGOTHERRECEIVED ;
output L0STATSCFGOTHERTRANSMITTED ;
output L0STATSCFGRECEIVED ;
output L0STATSCFGTRANSMITTED ;
output L0STATSDLLPRECEIVED ;
output L0STATSDLLPTRANSMITTED ;
output L0STATSOSRECEIVED ;
output L0STATSOSTRANSMITTED ;
output L0STATSTLPRECEIVED ;
output L0STATSTLPTRANSMITTED ;
output L0UNLOCKRECEIVED ;
output LLKRXEOFN ;
output LLKRXEOPN ;
output LLKRXSOFN ;
output LLKRXSOPN ;
output LLKRXSRCLASTREQN ;
output LLKRXSRCRDYN ;
output LLKTXCONFIGREADYN ;
output LLKTXDSTRDYN ;
output MEMSPACEENABLE ;
output MIMDLLBREN ;
output MIMDLLBWEN ;
output MIMRXBREN ;
output MIMRXBWEN ;
output MIMTXBREN ;
output MIMTXBWEN ;
output PARITYERRORRESPONSE ;
output PIPEDESKEWLANESL0 ;
output PIPEDESKEWLANESL1 ;
output PIPEDESKEWLANESL2 ;
output PIPEDESKEWLANESL3 ;
output PIPEDESKEWLANESL4 ;
output PIPEDESKEWLANESL5 ;
output PIPEDESKEWLANESL6 ;
output PIPEDESKEWLANESL7 ;
output PIPERESETL0 ;
output PIPERESETL1 ;
output PIPERESETL2 ;
output PIPERESETL3 ;
output PIPERESETL4 ;
output PIPERESETL5 ;
output PIPERESETL6 ;
output PIPERESETL7 ;
output PIPERXPOLARITYL0 ;
output PIPERXPOLARITYL1 ;
output PIPERXPOLARITYL2 ;
output PIPERXPOLARITYL3 ;
output PIPERXPOLARITYL4 ;
output PIPERXPOLARITYL5 ;
output PIPERXPOLARITYL6 ;
output PIPERXPOLARITYL7 ;
output PIPETXCOMPLIANCEL0 ;
output PIPETXCOMPLIANCEL1 ;
output PIPETXCOMPLIANCEL2 ;
output PIPETXCOMPLIANCEL3 ;
output PIPETXCOMPLIANCEL4 ;
output PIPETXCOMPLIANCEL5 ;
output PIPETXCOMPLIANCEL6 ;
output PIPETXCOMPLIANCEL7 ;
output PIPETXDATAKL0 ;
output PIPETXDATAKL1 ;
output PIPETXDATAKL2 ;
output PIPETXDATAKL3 ;
output PIPETXDATAKL4 ;
output PIPETXDATAKL5 ;
output PIPETXDATAKL6 ;
output PIPETXDATAKL7 ;
output PIPETXDETECTRXLOOPBACKL0 ;
output PIPETXDETECTRXLOOPBACKL1 ;
output PIPETXDETECTRXLOOPBACKL2 ;
output PIPETXDETECTRXLOOPBACKL3 ;
output PIPETXDETECTRXLOOPBACKL4 ;
output PIPETXDETECTRXLOOPBACKL5 ;
output PIPETXDETECTRXLOOPBACKL6 ;
output PIPETXDETECTRXLOOPBACKL7 ;
output PIPETXELECIDLEL0 ;
output PIPETXELECIDLEL1 ;
output PIPETXELECIDLEL2 ;
output PIPETXELECIDLEL3 ;
output PIPETXELECIDLEL4 ;
output PIPETXELECIDLEL5 ;
output PIPETXELECIDLEL6 ;
output PIPETXELECIDLEL7 ;
output SERRENABLE ;
output URREPORTINGENABLE ;
output [11:0] MGMTSTATSCREDIT ;
output [11:0] MIMDLLBRADD ;
output [11:0] MIMDLLBWADD ;
output [12:0] L0COMPLETERID ;
output [12:0] MIMRXBRADD ;
output [12:0] MIMRXBWADD ;
output [12:0] MIMTXBRADD ;
output [12:0] MIMTXBWADD ;
output [15:0] LLKRXPREFERREDTYPE ;
output [16:0] MGMTPSO ;
output [1:0] L0PWRSTATE0 ;
output [1:0] L0RXMACLINKERROR ;
output [1:0] LLKRXVALIDN ;
output [1:0] PIPEPOWERDOWNL0 ;
output [1:0] PIPEPOWERDOWNL1 ;
output [1:0] PIPEPOWERDOWNL2 ;
output [1:0] PIPEPOWERDOWNL3 ;
output [1:0] PIPEPOWERDOWNL4 ;
output [1:0] PIPEPOWERDOWNL5 ;
output [1:0] PIPEPOWERDOWNL6 ;
output [1:0] PIPEPOWERDOWNL7 ;
output [2:0] L0MULTIMSGEN0 ;
output [2:0] L0RXDLLPMTYPE ;
output [2:0] MAXPAYLOADSIZE ;
output [2:0] MAXREADREQUESTSIZE ;
output [31:0] MGMTRDATA ;
output [3:0] L0LTSSMSTATE ;
output [3:0] L0MACNEGOTIATEDLINKWIDTH ;
output [63:0] LLKRXDATA ;
output [63:0] MIMDLLBWDATA ;
output [63:0] MIMRXBWDATA ;
output [63:0] MIMTXBWDATA ;
output [6:0] L0DLLERRORVECTOR ;
output [7:0] L0DLLVCSTATUS ;
output [7:0] L0DLUPDOWN ;
output [7:0] LLKRXCHCOMPLETIONAVAILABLEN ;
output [7:0] LLKRXCHNONPOSTEDAVAILABLEN ;
output [7:0] LLKRXCHPOSTEDAVAILABLEN ;
output [7:0] LLKTCSTATUS ;
output [7:0] LLKTXCHCOMPLETIONREADYN ;
output [7:0] LLKTXCHNONPOSTEDREADYN ;
output [7:0] LLKTXCHPOSTEDREADYN ;
output [7:0] PIPETXDATAL0 ;
output [7:0] PIPETXDATAL1 ;
output [7:0] PIPETXDATAL2 ;
output [7:0] PIPETXDATAL3 ;
output [7:0] PIPETXDATAL4 ;
output [7:0] PIPETXDATAL5 ;
output [7:0] PIPETXDATAL6 ;
output [7:0] PIPETXDATAL7 ;
output [9:0] LLKTXCHANSPACE ;
parameter BAR0EXIST = "TRUE";
parameter BAR0PREFETCHABLE = "TRUE";
parameter BAR1EXIST = "FALSE";
parameter BAR1PREFETCHABLE = "FALSE";
parameter BAR2EXIST = "FALSE";
parameter BAR2PREFETCHABLE = "FALSE";
parameter BAR3EXIST = "FALSE";
parameter BAR3PREFETCHABLE = "FALSE";
parameter BAR4EXIST = "FALSE";
parameter BAR4PREFETCHABLE = "FALSE";
parameter BAR5EXIST = "FALSE";
parameter BAR5PREFETCHABLE = "FALSE";
parameter CLKDIVIDED = "FALSE";
parameter INFINITECOMPLETIONS = "TRUE";
parameter LINKSTATUSSLOTCLOCKCONFIG = "FALSE";
parameter PBCAPABILITYSYSTEMALLOCATED = "FALSE";
parameter PMCAPABILITYD1SUPPORT = "FALSE";
parameter PMCAPABILITYD2SUPPORT = "FALSE";
parameter PMCAPABILITYDSI = "TRUE";
parameter RESETMODE = "FALSE";
parameter [10:0] VC0TOTALCREDITSCD = 11'h0;
parameter [10:0] VC0TOTALCREDITSPD = 11'h34;
parameter [10:0] VC1TOTALCREDITSCD = 11'h0;
parameter [10:0] VC1TOTALCREDITSPD = 11'h0;
parameter [11:0] AERBASEPTR = 12'h110;
parameter [11:0] AERCAPABILITYNEXTPTR = 12'h138;
parameter [11:0] DSNBASEPTR = 12'h148;
parameter [11:0] DSNCAPABILITYNEXTPTR = 12'h154;
parameter [11:0] MSIBASEPTR = 12'h48;
parameter [11:0] PBBASEPTR = 12'h138;
parameter [11:0] PBCAPABILITYNEXTPTR = 12'h148;
parameter [11:0] PMBASEPTR = 12'h40;
parameter [11:0] RETRYRAMSIZE = 12'h9;
parameter [11:0] VCBASEPTR = 12'h154;
parameter [11:0] VCCAPABILITYNEXTPTR = 12'h0;
parameter [12:0] VC0RXFIFOBASEC = 13'h98;
parameter [12:0] VC0RXFIFOBASENP = 13'h80;
parameter [12:0] VC0RXFIFOBASEP = 13'h0;
parameter [12:0] VC0RXFIFOLIMITC = 13'h117;
parameter [12:0] VC0RXFIFOLIMITNP = 13'h97;
parameter [12:0] VC0RXFIFOLIMITP = 13'h7f;
parameter [12:0] VC0TXFIFOBASEC = 13'h98;
parameter [12:0] VC0TXFIFOBASENP = 13'h80;
parameter [12:0] VC0TXFIFOBASEP = 13'h0;
parameter [12:0] VC0TXFIFOLIMITC = 13'h117;
parameter [12:0] VC0TXFIFOLIMITNP = 13'h97;
parameter [12:0] VC0TXFIFOLIMITP = 13'h7f;
parameter [12:0] VC1RXFIFOBASEC = 13'h118;
parameter [12:0] VC1RXFIFOBASENP = 13'h118;
parameter [12:0] VC1RXFIFOBASEP = 13'h118;
parameter [12:0] VC1RXFIFOLIMITC = 13'h118;
parameter [12:0] VC1RXFIFOLIMITNP = 13'h118;
parameter [12:0] VC1RXFIFOLIMITP = 13'h118;
parameter [12:0] VC1TXFIFOBASEC = 13'h118;
parameter [12:0] VC1TXFIFOBASENP = 13'h118;
parameter [12:0] VC1TXFIFOBASEP = 13'h118;
parameter [12:0] VC1TXFIFOLIMITC = 13'h118;
parameter [12:0] VC1TXFIFOLIMITNP = 13'h118;
parameter [12:0] VC1TXFIFOLIMITP = 13'h118;
parameter [15:0] DEVICEID = 16'h5050;
parameter [15:0] SUBSYSTEMID = 16'h5050;
parameter [15:0] SUBSYSTEMVENDORID = 16'h10EE;
parameter [15:0] VENDORID = 16'h10EE;
parameter [1:0] LINKCAPABILITYASPMSUPPORT = 2'h1;
parameter [1:0] PBCAPABILITYDW0DATASCALE = 2'h0;
parameter [1:0] PBCAPABILITYDW0PMSTATE = 2'h0;
parameter [1:0] PBCAPABILITYDW1DATASCALE = 2'h0;
parameter [1:0] PBCAPABILITYDW1PMSTATE = 2'h0;
parameter [1:0] PBCAPABILITYDW2DATASCALE = 2'h0;
parameter [1:0] PBCAPABILITYDW2PMSTATE = 2'h0;
parameter [1:0] PBCAPABILITYDW3DATASCALE = 2'h0;
parameter [1:0] PBCAPABILITYDW3PMSTATE = 2'h0;
parameter [23:0] CLASSCODE = 24'h058000;
parameter [2:0] DEVICECAPABILITYENDPOINTL0SLATENCY = 3'h0;
parameter [2:0] DEVICECAPABILITYENDPOINTL1LATENCY = 3'h0;
parameter [2:0] MSICAPABILITYMULTIMSGCAP = 3'h0;
parameter [2:0] PBCAPABILITYDW0PMSUBSTATE = 3'h0;
parameter [2:0] PBCAPABILITYDW0POWERRAIL = 3'h0;
parameter [2:0] PBCAPABILITYDW0TYPE = 3'h0;
parameter [2:0] PBCAPABILITYDW1PMSUBSTATE = 3'h0;
parameter [2:0] PBCAPABILITYDW1POWERRAIL = 3'h0;
parameter [2:0] PBCAPABILITYDW1TYPE = 3'h0;
parameter [2:0] PBCAPABILITYDW2PMSUBSTATE = 3'h0;
parameter [2:0] PBCAPABILITYDW2POWERRAIL = 3'h0;
parameter [2:0] PBCAPABILITYDW2TYPE = 3'h0;
parameter [2:0] PBCAPABILITYDW3PMSUBSTATE = 3'h0;
parameter [2:0] PBCAPABILITYDW3POWERRAIL = 3'h0;
parameter [2:0] PBCAPABILITYDW3TYPE = 3'h0;
parameter [2:0] PMCAPABILITYAUXCURRENT = 3'h0;
parameter [2:0] PORTVCCAPABILITYEXTENDEDVCCOUNT = 3'h0;
parameter [31:0] CARDBUSCISPOINTER = 32'h0;
parameter [3:0] XPDEVICEPORTTYPE = 4'h0;
parameter [4:0] PMCAPABILITYPMESUPPORT = 5'h0;
parameter [5:0] BAR0MASKWIDTH = 6'h14;
parameter [5:0] BAR1MASKWIDTH = 6'h0;
parameter [5:0] BAR2MASKWIDTH = 6'h0;
parameter [5:0] BAR3MASKWIDTH = 6'h0;
parameter [5:0] BAR4MASKWIDTH = 6'h0;
parameter [5:0] BAR5MASKWIDTH = 6'h0;
parameter [5:0] LINKCAPABILITYMAXLINKWIDTH = 6'h01;
parameter [63:0] DEVICESERIALNUMBER = 64'hE000000001000A35;
parameter [6:0] VC0TOTALCREDITSCH = 7'h0;
parameter [6:0] VC0TOTALCREDITSNPH = 7'h08;
parameter [6:0] VC0TOTALCREDITSPH = 7'h08;
parameter [6:0] VC1TOTALCREDITSCH = 7'h0;
parameter [6:0] VC1TOTALCREDITSNPH = 7'h0;
parameter [6:0] VC1TOTALCREDITSPH = 7'h0;
parameter [7:0] ACTIVELANESIN = 8'h1;
parameter [7:0] CAPABILITIESPOINTER = 8'h40;
parameter [7:0] INTERRUPTPIN = 8'h0;
parameter [7:0] MSICAPABILITYNEXTPTR = 8'h60;
parameter [7:0] PBCAPABILITYDW0BASEPOWER = 8'h0;
parameter [7:0] PBCAPABILITYDW1BASEPOWER = 8'h0;
parameter [7:0] PBCAPABILITYDW2BASEPOWER = 8'h0;
parameter [7:0] PBCAPABILITYDW3BASEPOWER = 8'h0;
parameter [7:0] PCIECAPABILITYNEXTPTR = 8'h0;
parameter [7:0] PMCAPABILITYNEXTPTR = 8'h60;
parameter [7:0] PMDATA0 = 8'h0;
parameter [7:0] PMDATA1 = 8'h0;
parameter [7:0] PMDATA2 = 8'h0;
parameter [7:0] PMDATA3 = 8'h0;
parameter [7:0] PMDATA4 = 8'h0;
parameter [7:0] PMDATA5 = 8'h0;
parameter [7:0] PMDATA6 = 8'h0;
parameter [7:0] PMDATA7 = 8'h0;
parameter [7:0] PORTVCCAPABILITYVCARBCAP = 8'h0;
parameter [7:0] PORTVCCAPABILITYVCARBTABLEOFFSET = 8'h0;
parameter [7:0] REVISIONID = 8'h0;
parameter [7:0] XPBASEPTR = 8'h60;
parameter BAR0ADDRWIDTH = 0;
parameter BAR0IOMEMN = 0;
parameter BAR1ADDRWIDTH = 0;
parameter BAR1IOMEMN = 0;
parameter BAR2ADDRWIDTH = 0;
parameter BAR2IOMEMN = 0;
parameter BAR3ADDRWIDTH = 0;
parameter BAR3IOMEMN = 0;
parameter BAR4ADDRWIDTH = 0;
parameter BAR4IOMEMN = 0;
parameter BAR5IOMEMN = 0;
parameter L0SEXITLATENCY = 7;
parameter L0SEXITLATENCYCOMCLK = 7;
parameter L1EXITLATENCY = 7;
parameter L1EXITLATENCYCOMCLK = 7;
parameter LOWPRIORITYVCCOUNT = 0;
parameter PMDATASCALE0 = 0;
parameter PMDATASCALE1 = 0;
parameter PMDATASCALE2 = 0;
parameter PMDATASCALE3 = 0;
parameter PMDATASCALE4 = 0;
parameter PMDATASCALE5 = 0;
parameter PMDATASCALE6 = 0;
parameter PMDATASCALE7 = 0;
parameter RETRYRAMREADLATENCY = 3;
parameter RETRYRAMWRITELATENCY = 1;
parameter TLRAMREADLATENCY = 3;
parameter TLRAMWRITELATENCY = 1;
parameter TXTSNFTS = 255;
parameter TXTSNFTSCOMCLK = 255;
parameter XPMAXPAYLOAD = 0;
endmodule
//#### END MODULE DEFINITION FOR: PCIE_EP ####

//#### BEGIN MODULE DEFINITION FOR :PCIE_INTERNAL_1_1 ###
module PCIE_INTERNAL_1_1 (
	BUSMASTERENABLE,
	CRMDOHOTRESETN,
	CRMPWRSOFTRESETN,
	CRMRXHOTRESETN,
	DLLTXPMDLLPOUTSTANDING,
	INTERRUPTDISABLE,
	IOSPACEENABLE,
	L0ASAUTONOMOUSINITCOMPLETED,
	L0ATTENTIONINDICATORCONTROL,
	L0CFGLOOPBACKACK,
	L0COMPLETERID,
	L0CORRERRMSGRCVD,
	L0DLLASRXSTATE,
	L0DLLASTXSTATE,
	L0DLLERRORVECTOR,
	L0DLLRXACKOUTSTANDING,
	L0DLLTXNONFCOUTSTANDING,
	L0DLLTXOUTSTANDING,
	L0DLLVCSTATUS,
	L0DLUPDOWN,
	L0ERRMSGREQID,
	L0FATALERRMSGRCVD,
	L0FIRSTCFGWRITEOCCURRED,
	L0FWDCORRERROUT,
	L0FWDFATALERROUT,
	L0FWDNONFATALERROUT,
	L0LTSSMSTATE,
	L0MACENTEREDL0,
	L0MACLINKTRAINING,
	L0MACLINKUP,
	L0MACNEGOTIATEDLINKWIDTH,
	L0MACNEWSTATEACK,
	L0MACRXL0SSTATE,
	L0MACUPSTREAMDOWNSTREAM,
	L0MCFOUND,
	L0MSIENABLE0,
	L0MULTIMSGEN0,
	L0NONFATALERRMSGRCVD,
	L0PMEACK,
	L0PMEEN,
	L0PMEREQOUT,
	L0POWERCONTROLLERCONTROL,
	L0POWERINDICATORCONTROL,
	L0PWRINHIBITTRANSFERS,
	L0PWRL1STATE,
	L0PWRL23READYDEVICE,
	L0PWRL23READYSTATE,
	L0PWRSTATE0,
	L0PWRTURNOFFREQ,
	L0PWRTXL0SSTATE,
	L0RECEIVEDASSERTINTALEGACYINT,
	L0RECEIVEDASSERTINTBLEGACYINT,
	L0RECEIVEDASSERTINTCLEGACYINT,
	L0RECEIVEDASSERTINTDLEGACYINT,
	L0RECEIVEDDEASSERTINTALEGACYINT,
	L0RECEIVEDDEASSERTINTBLEGACYINT,
	L0RECEIVEDDEASSERTINTCLEGACYINT,
	L0RECEIVEDDEASSERTINTDLEGACYINT,
	L0RXBEACON,
	L0RXDLLFCCMPLMCCRED,
	L0RXDLLFCCMPLMCUPDATE,
	L0RXDLLFCNPOSTBYPCRED,
	L0RXDLLFCNPOSTBYPUPDATE,
	L0RXDLLFCPOSTORDCRED,
	L0RXDLLFCPOSTORDUPDATE,
	L0RXDLLPM,
	L0RXDLLPMTYPE,
	L0RXDLLSBFCDATA,
	L0RXDLLSBFCUPDATE,
	L0RXDLLTLPECRCOK,
	L0RXDLLTLPEND,
	L0RXMACLINKERROR,
	L0STATSCFGOTHERRECEIVED,
	L0STATSCFGOTHERTRANSMITTED,
	L0STATSCFGRECEIVED,
	L0STATSCFGTRANSMITTED,
	L0STATSDLLPRECEIVED,
	L0STATSDLLPTRANSMITTED,
	L0STATSOSRECEIVED,
	L0STATSOSTRANSMITTED,
	L0STATSTLPRECEIVED,
	L0STATSTLPTRANSMITTED,
	L0TOGGLEELECTROMECHANICALINTERLOCK,
	L0TRANSFORMEDVC,
	L0TXDLLFCCMPLMCUPDATED,
	L0TXDLLFCNPOSTBYPUPDATED,
	L0TXDLLFCPOSTORDUPDATED,
	L0TXDLLPMUPDATED,
	L0TXDLLSBFCUPDATED,
	L0UCBYPFOUND,
	L0UCORDFOUND,
	L0UNLOCKRECEIVED,
	LLKRX4DWHEADERN,
	LLKRXCHCOMPLETIONAVAILABLEN,
	LLKRXCHCOMPLETIONPARTIALN,
	LLKRXCHCONFIGAVAILABLEN,
	LLKRXCHCONFIGPARTIALN,
	LLKRXCHNONPOSTEDAVAILABLEN,
	LLKRXCHNONPOSTEDPARTIALN,
	LLKRXCHPOSTEDAVAILABLEN,
	LLKRXCHPOSTEDPARTIALN,
	LLKRXDATA,
	LLKRXECRCBADN,
	LLKRXEOFN,
	LLKRXEOPN,
	LLKRXPREFERREDTYPE,
	LLKRXSOFN,
	LLKRXSOPN,
	LLKRXSRCDSCN,
	LLKRXSRCLASTREQN,
	LLKRXSRCRDYN,
	LLKRXVALIDN,
	LLKTCSTATUS,
	LLKTXCHANSPACE,
	LLKTXCHCOMPLETIONREADYN,
	LLKTXCHNONPOSTEDREADYN,
	LLKTXCHPOSTEDREADYN,
	LLKTXCONFIGREADYN,
	LLKTXDSTRDYN,
	MAXPAYLOADSIZE,
	MAXREADREQUESTSIZE,
	MEMSPACEENABLE,
	MGMTPSO,
	MGMTRDATA,
	MGMTSTATSCREDIT,
	MIMDLLBRADD,
	MIMDLLBREN,
	MIMDLLBWADD,
	MIMDLLBWDATA,
	MIMDLLBWEN,
	MIMRXBRADD,
	MIMRXBREN,
	MIMRXBWADD,
	MIMRXBWDATA,
	MIMRXBWEN,
	MIMTXBRADD,
	MIMTXBREN,
	MIMTXBWADD,
	MIMTXBWDATA,
	MIMTXBWEN,
	PARITYERRORRESPONSE,
	PIPEDESKEWLANESL0,
	PIPEDESKEWLANESL1,
	PIPEDESKEWLANESL2,
	PIPEDESKEWLANESL3,
	PIPEDESKEWLANESL4,
	PIPEDESKEWLANESL5,
	PIPEDESKEWLANESL6,
	PIPEDESKEWLANESL7,
	PIPEPOWERDOWNL0,
	PIPEPOWERDOWNL1,
	PIPEPOWERDOWNL2,
	PIPEPOWERDOWNL3,
	PIPEPOWERDOWNL4,
	PIPEPOWERDOWNL5,
	PIPEPOWERDOWNL6,
	PIPEPOWERDOWNL7,
	PIPERESETL0,
	PIPERESETL1,
	PIPERESETL2,
	PIPERESETL3,
	PIPERESETL4,
	PIPERESETL5,
	PIPERESETL6,
	PIPERESETL7,
	PIPERXPOLARITYL0,
	PIPERXPOLARITYL1,
	PIPERXPOLARITYL2,
	PIPERXPOLARITYL3,
	PIPERXPOLARITYL4,
	PIPERXPOLARITYL5,
	PIPERXPOLARITYL6,
	PIPERXPOLARITYL7,
	PIPETXCOMPLIANCEL0,
	PIPETXCOMPLIANCEL1,
	PIPETXCOMPLIANCEL2,
	PIPETXCOMPLIANCEL3,
	PIPETXCOMPLIANCEL4,
	PIPETXCOMPLIANCEL5,
	PIPETXCOMPLIANCEL6,
	PIPETXCOMPLIANCEL7,
	PIPETXDATAKL0,
	PIPETXDATAKL1,
	PIPETXDATAKL2,
	PIPETXDATAKL3,
	PIPETXDATAKL4,
	PIPETXDATAKL5,
	PIPETXDATAKL6,
	PIPETXDATAKL7,
	PIPETXDATAL0,
	PIPETXDATAL1,
	PIPETXDATAL2,
	PIPETXDATAL3,
	PIPETXDATAL4,
	PIPETXDATAL5,
	PIPETXDATAL6,
	PIPETXDATAL7,
	PIPETXDETECTRXLOOPBACKL0,
	PIPETXDETECTRXLOOPBACKL1,
	PIPETXDETECTRXLOOPBACKL2,
	PIPETXDETECTRXLOOPBACKL3,
	PIPETXDETECTRXLOOPBACKL4,
	PIPETXDETECTRXLOOPBACKL5,
	PIPETXDETECTRXLOOPBACKL6,
	PIPETXDETECTRXLOOPBACKL7,
	PIPETXELECIDLEL0,
	PIPETXELECIDLEL1,
	PIPETXELECIDLEL2,
	PIPETXELECIDLEL3,
	PIPETXELECIDLEL4,
	PIPETXELECIDLEL5,
	PIPETXELECIDLEL6,
	PIPETXELECIDLEL7,
	SERRENABLE,
	URREPORTINGENABLE,

	AUXPOWER,
	CFGNEGOTIATEDLINKWIDTH,
	COMPLIANCEAVOID,
	CRMCFGBRIDGEHOTRESET,
	CRMCORECLK,
	CRMCORECLKDLO,
	CRMCORECLKRXO,
	CRMCORECLKTXO,
	CRMLINKRSTN,
	CRMMACRSTN,
	CRMMGMTRSTN,
	CRMNVRSTN,
	CRMTXHOTRESETN,
	CRMURSTN,
	CRMUSERCFGRSTN,
	CRMUSERCLK,
	CRMUSERCLKRXO,
	CRMUSERCLKTXO,
	CROSSLINKSEED,
	L0ACKNAKTIMERADJUSTMENT,
	L0ALLDOWNPORTSINL1,
	L0ALLDOWNRXPORTSINL0S,
	L0ASE,
	L0ASPORTCOUNT,
	L0ASTURNPOOLBITSCONSUMED,
	L0ATTENTIONBUTTONPRESSED,
	L0CFGASSPANTREEOWNEDSTATE,
	L0CFGASSTATECHANGECMD,
	L0CFGDISABLESCRAMBLE,
	L0CFGEXTENDEDSYNC,
	L0CFGL0SENTRYENABLE,
	L0CFGL0SENTRYSUP,
	L0CFGL0SEXITLAT,
	L0CFGLINKDISABLE,
	L0CFGLOOPBACKMASTER,
	L0CFGNEGOTIATEDMAXP,
	L0CFGVCENABLE,
	L0CFGVCID,
	L0DLLHOLDLINKUP,
	L0ELECTROMECHANICALINTERLOCKENGAGED,
	L0FWDASSERTINTALEGACYINT,
	L0FWDASSERTINTBLEGACYINT,
	L0FWDASSERTINTCLEGACYINT,
	L0FWDASSERTINTDLEGACYINT,
	L0FWDCORRERRIN,
	L0FWDDEASSERTINTALEGACYINT,
	L0FWDDEASSERTINTBLEGACYINT,
	L0FWDDEASSERTINTCLEGACYINT,
	L0FWDDEASSERTINTDLEGACYINT,
	L0FWDFATALERRIN,
	L0FWDNONFATALERRIN,
	L0LEGACYINTFUNCT0,
	L0MRLSENSORCLOSEDN,
	L0MSIREQUEST0,
	L0PACKETHEADERFROMUSER,
	L0PMEREQIN,
	L0PORTNUMBER,
	L0POWERFAULTDETECTED,
	L0PRESENCEDETECTSLOTEMPTYN,
	L0PWRNEWSTATEREQ,
	L0PWRNEXTLINKSTATE,
	L0REPLAYTIMERADJUSTMENT,
	L0ROOTTURNOFFREQ,
	L0RXTLTLPNONINITIALIZEDVC,
	L0SENDUNLOCKMESSAGE,
	L0SETCOMPLETERABORTERROR,
	L0SETCOMPLETIONTIMEOUTCORRERROR,
	L0SETCOMPLETIONTIMEOUTUNCORRERROR,
	L0SETDETECTEDCORRERROR,
	L0SETDETECTEDFATALERROR,
	L0SETDETECTEDNONFATALERROR,
	L0SETLINKDETECTEDPARITYERROR,
	L0SETLINKMASTERDATAPARITY,
	L0SETLINKRECEIVEDMASTERABORT,
	L0SETLINKRECEIVEDTARGETABORT,
	L0SETLINKSIGNALLEDTARGETABORT,
	L0SETLINKSYSTEMERROR,
	L0SETUNEXPECTEDCOMPLETIONCORRERROR,
	L0SETUNEXPECTEDCOMPLETIONUNCORRERROR,
	L0SETUNSUPPORTEDREQUESTNONPOSTEDERROR,
	L0SETUNSUPPORTEDREQUESTOTHERERROR,
	L0SETUSERDETECTEDPARITYERROR,
	L0SETUSERMASTERDATAPARITY,
	L0SETUSERRECEIVEDMASTERABORT,
	L0SETUSERRECEIVEDTARGETABORT,
	L0SETUSERSIGNALLEDTARGETABORT,
	L0SETUSERSYSTEMERROR,
	L0TLASFCCREDSTARVATION,
	L0TLLINKRETRAIN,
	L0TRANSACTIONSPENDING,
	L0TXBEACON,
	L0TXCFGPM,
	L0TXCFGPMTYPE,
	L0TXTLFCCMPLMCCRED,
	L0TXTLFCCMPLMCUPDATE,
	L0TXTLFCNPOSTBYPCRED,
	L0TXTLFCNPOSTBYPUPDATE,
	L0TXTLFCPOSTORDCRED,
	L0TXTLFCPOSTORDUPDATE,
	L0TXTLSBFCDATA,
	L0TXTLSBFCUPDATE,
	L0TXTLTLPDATA,
	L0TXTLTLPEDB,
	L0TXTLTLPENABLE,
	L0TXTLTLPEND,
	L0TXTLTLPLATENCY,
	L0TXTLTLPREQ,
	L0TXTLTLPREQEND,
	L0TXTLTLPWIDTH,
	L0UPSTREAMRXPORTINL0S,
	L0VC0PREVIEWEXPAND,
	L0WAKEN,
	LLKRXCHFIFO,
	LLKRXCHTC,
	LLKRXDSTCONTREQN,
	LLKRXDSTREQN,
	LLKTX4DWHEADERN,
	LLKTXCHFIFO,
	LLKTXCHTC,
	LLKTXCOMPLETEN,
	LLKTXCREATEECRCN,
	LLKTXDATA,
	LLKTXENABLEN,
	LLKTXEOFN,
	LLKTXEOPN,
	LLKTXSOFN,
	LLKTXSOPN,
	LLKTXSRCDSCN,
	LLKTXSRCRDYN,
	MAINPOWER,
	MGMTADDR,
	MGMTBWREN,
	MGMTRDEN,
	MGMTSTATSCREDITSEL,
	MGMTWDATA,
	MGMTWREN,
	MIMDLLBRDATA,
	MIMRXBRDATA,
	MIMTXBRDATA,
	PIPEPHYSTATUSL0,
	PIPEPHYSTATUSL1,
	PIPEPHYSTATUSL2,
	PIPEPHYSTATUSL3,
	PIPEPHYSTATUSL4,
	PIPEPHYSTATUSL5,
	PIPEPHYSTATUSL6,
	PIPEPHYSTATUSL7,
	PIPERXCHANISALIGNEDL0,
	PIPERXCHANISALIGNEDL1,
	PIPERXCHANISALIGNEDL2,
	PIPERXCHANISALIGNEDL3,
	PIPERXCHANISALIGNEDL4,
	PIPERXCHANISALIGNEDL5,
	PIPERXCHANISALIGNEDL6,
	PIPERXCHANISALIGNEDL7,
	PIPERXDATAKL0,
	PIPERXDATAKL1,
	PIPERXDATAKL2,
	PIPERXDATAKL3,
	PIPERXDATAKL4,
	PIPERXDATAKL5,
	PIPERXDATAKL6,
	PIPERXDATAKL7,
	PIPERXDATAL0,
	PIPERXDATAL1,
	PIPERXDATAL2,
	PIPERXDATAL3,
	PIPERXDATAL4,
	PIPERXDATAL5,
	PIPERXDATAL6,
	PIPERXDATAL7,
	PIPERXELECIDLEL0,
	PIPERXELECIDLEL1,
	PIPERXELECIDLEL2,
	PIPERXELECIDLEL3,
	PIPERXELECIDLEL4,
	PIPERXELECIDLEL5,
	PIPERXELECIDLEL6,
	PIPERXELECIDLEL7,
	PIPERXSTATUSL0,
	PIPERXSTATUSL1,
	PIPERXSTATUSL2,
	PIPERXSTATUSL3,
	PIPERXSTATUSL4,
	PIPERXSTATUSL5,
	PIPERXSTATUSL6,
	PIPERXSTATUSL7,
	PIPERXVALIDL0,
	PIPERXVALIDL1,
	PIPERXVALIDL2,
	PIPERXVALIDL3,
	PIPERXVALIDL4,
	PIPERXVALIDL5,
	PIPERXVALIDL6,
	PIPERXVALIDL7

) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input AUXPOWER ;
input COMPLIANCEAVOID ;
input CRMCFGBRIDGEHOTRESET ;
input CRMCORECLK ;
input CRMCORECLKDLO ;
input CRMCORECLKRXO ;
input CRMCORECLKTXO ;
input CRMLINKRSTN ;
input CRMMACRSTN ;
input CRMMGMTRSTN ;
input CRMNVRSTN ;
input CRMTXHOTRESETN ;
input CRMURSTN ;
input CRMUSERCFGRSTN ;
input CRMUSERCLK ;
input CRMUSERCLKRXO ;
input CRMUSERCLKTXO ;
input CROSSLINKSEED ;
input L0ALLDOWNPORTSINL1 ;
input L0ALLDOWNRXPORTSINL0S ;
input L0ASE ;
input L0ATTENTIONBUTTONPRESSED ;
input L0CFGASSPANTREEOWNEDSTATE ;
input L0CFGDISABLESCRAMBLE ;
input L0CFGEXTENDEDSYNC ;
input L0CFGL0SENTRYENABLE ;
input L0CFGL0SENTRYSUP ;
input L0CFGLINKDISABLE ;
input L0CFGLOOPBACKMASTER ;
input L0DLLHOLDLINKUP ;
input L0ELECTROMECHANICALINTERLOCKENGAGED ;
input L0FWDASSERTINTALEGACYINT ;
input L0FWDASSERTINTBLEGACYINT ;
input L0FWDASSERTINTCLEGACYINT ;
input L0FWDASSERTINTDLEGACYINT ;
input L0FWDCORRERRIN ;
input L0FWDDEASSERTINTALEGACYINT ;
input L0FWDDEASSERTINTBLEGACYINT ;
input L0FWDDEASSERTINTCLEGACYINT ;
input L0FWDDEASSERTINTDLEGACYINT ;
input L0FWDFATALERRIN ;
input L0FWDNONFATALERRIN ;
input L0LEGACYINTFUNCT0 ;
input L0MRLSENSORCLOSEDN ;
input L0PMEREQIN ;
input L0POWERFAULTDETECTED ;
input L0PRESENCEDETECTSLOTEMPTYN ;
input L0PWRNEWSTATEREQ ;
input L0ROOTTURNOFFREQ ;
input L0SENDUNLOCKMESSAGE ;
input L0SETCOMPLETERABORTERROR ;
input L0SETCOMPLETIONTIMEOUTCORRERROR ;
input L0SETCOMPLETIONTIMEOUTUNCORRERROR ;
input L0SETDETECTEDCORRERROR ;
input L0SETDETECTEDFATALERROR ;
input L0SETDETECTEDNONFATALERROR ;
input L0SETLINKDETECTEDPARITYERROR ;
input L0SETLINKMASTERDATAPARITY ;
input L0SETLINKRECEIVEDMASTERABORT ;
input L0SETLINKRECEIVEDTARGETABORT ;
input L0SETLINKSIGNALLEDTARGETABORT ;
input L0SETLINKSYSTEMERROR ;
input L0SETUNEXPECTEDCOMPLETIONCORRERROR ;
input L0SETUNEXPECTEDCOMPLETIONUNCORRERROR ;
input L0SETUNSUPPORTEDREQUESTNONPOSTEDERROR ;
input L0SETUNSUPPORTEDREQUESTOTHERERROR ;
input L0SETUSERDETECTEDPARITYERROR ;
input L0SETUSERMASTERDATAPARITY ;
input L0SETUSERRECEIVEDMASTERABORT ;
input L0SETUSERRECEIVEDTARGETABORT ;
input L0SETUSERSIGNALLEDTARGETABORT ;
input L0SETUSERSYSTEMERROR ;
input L0TLASFCCREDSTARVATION ;
input L0TLLINKRETRAIN ;
input L0TRANSACTIONSPENDING ;
input L0TXBEACON ;
input L0TXCFGPM ;
input L0TXTLSBFCUPDATE ;
input L0TXTLTLPEDB ;
input L0TXTLTLPREQ ;
input L0TXTLTLPREQEND ;
input L0TXTLTLPWIDTH ;
input L0UPSTREAMRXPORTINL0S ;
input L0VC0PREVIEWEXPAND ;
input L0WAKEN ;
input LLKRXDSTCONTREQN ;
input LLKRXDSTREQN ;
input LLKTX4DWHEADERN ;
input LLKTXCOMPLETEN ;
input LLKTXCREATEECRCN ;
input LLKTXEOFN ;
input LLKTXEOPN ;
input LLKTXSOFN ;
input LLKTXSOPN ;
input LLKTXSRCDSCN ;
input LLKTXSRCRDYN ;
input MAINPOWER ;
input MGMTRDEN ;
input MGMTWREN ;
input PIPEPHYSTATUSL0 ;
input PIPEPHYSTATUSL1 ;
input PIPEPHYSTATUSL2 ;
input PIPEPHYSTATUSL3 ;
input PIPEPHYSTATUSL4 ;
input PIPEPHYSTATUSL5 ;
input PIPEPHYSTATUSL6 ;
input PIPEPHYSTATUSL7 ;
input PIPERXCHANISALIGNEDL0 ;
input PIPERXCHANISALIGNEDL1 ;
input PIPERXCHANISALIGNEDL2 ;
input PIPERXCHANISALIGNEDL3 ;
input PIPERXCHANISALIGNEDL4 ;
input PIPERXCHANISALIGNEDL5 ;
input PIPERXCHANISALIGNEDL6 ;
input PIPERXCHANISALIGNEDL7 ;
input PIPERXDATAKL0 ;
input PIPERXDATAKL1 ;
input PIPERXDATAKL2 ;
input PIPERXDATAKL3 ;
input PIPERXDATAKL4 ;
input PIPERXDATAKL5 ;
input PIPERXDATAKL6 ;
input PIPERXDATAKL7 ;
input PIPERXELECIDLEL0 ;
input PIPERXELECIDLEL1 ;
input PIPERXELECIDLEL2 ;
input PIPERXELECIDLEL3 ;
input PIPERXELECIDLEL4 ;
input PIPERXELECIDLEL5 ;
input PIPERXELECIDLEL6 ;
input PIPERXELECIDLEL7 ;
input PIPERXVALIDL0 ;
input PIPERXVALIDL1 ;
input PIPERXVALIDL2 ;
input PIPERXVALIDL3 ;
input PIPERXVALIDL4 ;
input PIPERXVALIDL5 ;
input PIPERXVALIDL6 ;
input PIPERXVALIDL7 ;
input [10:0] MGMTADDR ;
input [11:0] L0ACKNAKTIMERADJUSTMENT ;
input [11:0] L0REPLAYTIMERADJUSTMENT ;
input [127:0] L0PACKETHEADERFROMUSER ;
input [159:0] L0TXTLFCCMPLMCCRED ;
input [159:0] L0TXTLFCPOSTORDCRED ;
input [15:0] L0TXTLFCCMPLMCUPDATE ;
input [15:0] L0TXTLFCNPOSTBYPUPDATE ;
input [15:0] L0TXTLFCPOSTORDUPDATE ;
input [18:0] L0TXTLSBFCDATA ;
input [191:0] L0TXTLFCNPOSTBYPCRED ;
input [1:0] L0PWRNEXTLINKSTATE ;
input [1:0] L0TXTLTLPENABLE ;
input [1:0] L0TXTLTLPEND ;
input [1:0] LLKRXCHFIFO ;
input [1:0] LLKTXCHFIFO ;
input [1:0] LLKTXENABLEN ;
input [23:0] L0CFGVCID ;
input [2:0] L0ASTURNPOOLBITSCONSUMED ;
input [2:0] L0CFGL0SEXITLAT ;
input [2:0] L0CFGNEGOTIATEDMAXP ;
input [2:0] L0TXCFGPMTYPE ;
input [2:0] LLKRXCHTC ;
input [2:0] LLKTXCHTC ;
input [2:0] PIPERXSTATUSL0 ;
input [2:0] PIPERXSTATUSL1 ;
input [2:0] PIPERXSTATUSL2 ;
input [2:0] PIPERXSTATUSL3 ;
input [2:0] PIPERXSTATUSL4 ;
input [2:0] PIPERXSTATUSL5 ;
input [2:0] PIPERXSTATUSL6 ;
input [2:0] PIPERXSTATUSL7 ;
input [31:0] MGMTWDATA ;
input [3:0] L0CFGASSTATECHANGECMD ;
input [3:0] L0MSIREQUEST0 ;
input [3:0] L0TXTLTLPLATENCY ;
input [3:0] MGMTBWREN ;
input [5:0] CFGNEGOTIATEDLINKWIDTH ;
input [63:0] L0TXTLTLPDATA ;
input [63:0] LLKTXDATA ;
input [63:0] MIMDLLBRDATA ;
input [63:0] MIMRXBRDATA ;
input [63:0] MIMTXBRDATA ;
input [6:0] MGMTSTATSCREDITSEL ;
input [7:0] L0ASPORTCOUNT ;
input [7:0] L0CFGVCENABLE ;
input [7:0] L0PORTNUMBER ;
input [7:0] L0RXTLTLPNONINITIALIZEDVC ;
input [7:0] PIPERXDATAL0 ;
input [7:0] PIPERXDATAL1 ;
input [7:0] PIPERXDATAL2 ;
input [7:0] PIPERXDATAL3 ;
input [7:0] PIPERXDATAL4 ;
input [7:0] PIPERXDATAL5 ;
input [7:0] PIPERXDATAL6 ;
input [7:0] PIPERXDATAL7 ;
output BUSMASTERENABLE ;
output CRMDOHOTRESETN ;
output CRMPWRSOFTRESETN ;
output CRMRXHOTRESETN ;
output DLLTXPMDLLPOUTSTANDING ;
output INTERRUPTDISABLE ;
output IOSPACEENABLE ;
output L0ASAUTONOMOUSINITCOMPLETED ;
output L0CFGLOOPBACKACK ;
output L0CORRERRMSGRCVD ;
output L0DLLASTXSTATE ;
output L0DLLRXACKOUTSTANDING ;
output L0DLLTXNONFCOUTSTANDING ;
output L0DLLTXOUTSTANDING ;
output L0FATALERRMSGRCVD ;
output L0FIRSTCFGWRITEOCCURRED ;
output L0FWDCORRERROUT ;
output L0FWDFATALERROUT ;
output L0FWDNONFATALERROUT ;
output L0MACENTEREDL0 ;
output L0MACLINKTRAINING ;
output L0MACLINKUP ;
output L0MACNEWSTATEACK ;
output L0MACRXL0SSTATE ;
output L0MACUPSTREAMDOWNSTREAM ;
output L0MSIENABLE0 ;
output L0NONFATALERRMSGRCVD ;
output L0PMEACK ;
output L0PMEEN ;
output L0PMEREQOUT ;
output L0POWERCONTROLLERCONTROL ;
output L0PWRINHIBITTRANSFERS ;
output L0PWRL1STATE ;
output L0PWRL23READYDEVICE ;
output L0PWRL23READYSTATE ;
output L0PWRTURNOFFREQ ;
output L0PWRTXL0SSTATE ;
output L0RECEIVEDASSERTINTALEGACYINT ;
output L0RECEIVEDASSERTINTBLEGACYINT ;
output L0RECEIVEDASSERTINTCLEGACYINT ;
output L0RECEIVEDASSERTINTDLEGACYINT ;
output L0RECEIVEDDEASSERTINTALEGACYINT ;
output L0RECEIVEDDEASSERTINTBLEGACYINT ;
output L0RECEIVEDDEASSERTINTCLEGACYINT ;
output L0RECEIVEDDEASSERTINTDLEGACYINT ;
output L0RXBEACON ;
output L0RXDLLPM ;
output L0RXDLLSBFCUPDATE ;
output L0RXDLLTLPECRCOK ;
output L0STATSCFGOTHERRECEIVED ;
output L0STATSCFGOTHERTRANSMITTED ;
output L0STATSCFGRECEIVED ;
output L0STATSCFGTRANSMITTED ;
output L0STATSDLLPRECEIVED ;
output L0STATSDLLPTRANSMITTED ;
output L0STATSOSRECEIVED ;
output L0STATSOSTRANSMITTED ;
output L0STATSTLPRECEIVED ;
output L0STATSTLPTRANSMITTED ;
output L0TOGGLEELECTROMECHANICALINTERLOCK ;
output L0TXDLLPMUPDATED ;
output L0TXDLLSBFCUPDATED ;
output L0UNLOCKRECEIVED ;
output LLKRX4DWHEADERN ;
output LLKRXCHCONFIGAVAILABLEN ;
output LLKRXCHCONFIGPARTIALN ;
output LLKRXECRCBADN ;
output LLKRXEOFN ;
output LLKRXEOPN ;
output LLKRXSOFN ;
output LLKRXSOPN ;
output LLKRXSRCDSCN ;
output LLKRXSRCLASTREQN ;
output LLKRXSRCRDYN ;
output LLKTXCONFIGREADYN ;
output LLKTXDSTRDYN ;
output MEMSPACEENABLE ;
output MIMDLLBREN ;
output MIMDLLBWEN ;
output MIMRXBREN ;
output MIMRXBWEN ;
output MIMTXBREN ;
output MIMTXBWEN ;
output PARITYERRORRESPONSE ;
output PIPEDESKEWLANESL0 ;
output PIPEDESKEWLANESL1 ;
output PIPEDESKEWLANESL2 ;
output PIPEDESKEWLANESL3 ;
output PIPEDESKEWLANESL4 ;
output PIPEDESKEWLANESL5 ;
output PIPEDESKEWLANESL6 ;
output PIPEDESKEWLANESL7 ;
output PIPERESETL0 ;
output PIPERESETL1 ;
output PIPERESETL2 ;
output PIPERESETL3 ;
output PIPERESETL4 ;
output PIPERESETL5 ;
output PIPERESETL6 ;
output PIPERESETL7 ;
output PIPERXPOLARITYL0 ;
output PIPERXPOLARITYL1 ;
output PIPERXPOLARITYL2 ;
output PIPERXPOLARITYL3 ;
output PIPERXPOLARITYL4 ;
output PIPERXPOLARITYL5 ;
output PIPERXPOLARITYL6 ;
output PIPERXPOLARITYL7 ;
output PIPETXCOMPLIANCEL0 ;
output PIPETXCOMPLIANCEL1 ;
output PIPETXCOMPLIANCEL2 ;
output PIPETXCOMPLIANCEL3 ;
output PIPETXCOMPLIANCEL4 ;
output PIPETXCOMPLIANCEL5 ;
output PIPETXCOMPLIANCEL6 ;
output PIPETXCOMPLIANCEL7 ;
output PIPETXDATAKL0 ;
output PIPETXDATAKL1 ;
output PIPETXDATAKL2 ;
output PIPETXDATAKL3 ;
output PIPETXDATAKL4 ;
output PIPETXDATAKL5 ;
output PIPETXDATAKL6 ;
output PIPETXDATAKL7 ;
output PIPETXDETECTRXLOOPBACKL0 ;
output PIPETXDETECTRXLOOPBACKL1 ;
output PIPETXDETECTRXLOOPBACKL2 ;
output PIPETXDETECTRXLOOPBACKL3 ;
output PIPETXDETECTRXLOOPBACKL4 ;
output PIPETXDETECTRXLOOPBACKL5 ;
output PIPETXDETECTRXLOOPBACKL6 ;
output PIPETXDETECTRXLOOPBACKL7 ;
output PIPETXELECIDLEL0 ;
output PIPETXELECIDLEL1 ;
output PIPETXELECIDLEL2 ;
output PIPETXELECIDLEL3 ;
output PIPETXELECIDLEL4 ;
output PIPETXELECIDLEL5 ;
output PIPETXELECIDLEL6 ;
output PIPETXELECIDLEL7 ;
output SERRENABLE ;
output URREPORTINGENABLE ;
output [11:0] MGMTSTATSCREDIT ;
output [11:0] MIMDLLBRADD ;
output [11:0] MIMDLLBWADD ;
output [12:0] L0COMPLETERID ;
output [12:0] MIMRXBRADD ;
output [12:0] MIMRXBWADD ;
output [12:0] MIMTXBRADD ;
output [12:0] MIMTXBWADD ;
output [15:0] L0ERRMSGREQID ;
output [15:0] LLKRXPREFERREDTYPE ;
output [16:0] MGMTPSO ;
output [18:0] L0RXDLLSBFCDATA ;
output [19:0] L0RXDLLFCNPOSTBYPCRED ;
output [1:0] L0ATTENTIONINDICATORCONTROL ;
output [1:0] L0DLLASRXSTATE ;
output [1:0] L0POWERINDICATORCONTROL ;
output [1:0] L0PWRSTATE0 ;
output [1:0] L0RXDLLTLPEND ;
output [1:0] L0RXMACLINKERROR ;
output [1:0] LLKRXVALIDN ;
output [1:0] PIPEPOWERDOWNL0 ;
output [1:0] PIPEPOWERDOWNL1 ;
output [1:0] PIPEPOWERDOWNL2 ;
output [1:0] PIPEPOWERDOWNL3 ;
output [1:0] PIPEPOWERDOWNL4 ;
output [1:0] PIPEPOWERDOWNL5 ;
output [1:0] PIPEPOWERDOWNL6 ;
output [1:0] PIPEPOWERDOWNL7 ;
output [23:0] L0RXDLLFCCMPLMCCRED ;
output [23:0] L0RXDLLFCPOSTORDCRED ;
output [2:0] L0MCFOUND ;
output [2:0] L0MULTIMSGEN0 ;
output [2:0] L0RXDLLPMTYPE ;
output [2:0] L0TRANSFORMEDVC ;
output [2:0] MAXPAYLOADSIZE ;
output [2:0] MAXREADREQUESTSIZE ;
output [31:0] MGMTRDATA ;
output [3:0] L0LTSSMSTATE ;
output [3:0] L0MACNEGOTIATEDLINKWIDTH ;
output [3:0] L0UCBYPFOUND ;
output [3:0] L0UCORDFOUND ;
output [63:0] LLKRXDATA ;
output [63:0] MIMDLLBWDATA ;
output [63:0] MIMRXBWDATA ;
output [63:0] MIMTXBWDATA ;
output [6:0] L0DLLERRORVECTOR ;
output [7:0] L0DLLVCSTATUS ;
output [7:0] L0DLUPDOWN ;
output [7:0] L0RXDLLFCCMPLMCUPDATE ;
output [7:0] L0RXDLLFCNPOSTBYPUPDATE ;
output [7:0] L0RXDLLFCPOSTORDUPDATE ;
output [7:0] L0TXDLLFCCMPLMCUPDATED ;
output [7:0] L0TXDLLFCNPOSTBYPUPDATED ;
output [7:0] L0TXDLLFCPOSTORDUPDATED ;
output [7:0] LLKRXCHCOMPLETIONAVAILABLEN ;
output [7:0] LLKRXCHCOMPLETIONPARTIALN ;
output [7:0] LLKRXCHNONPOSTEDAVAILABLEN ;
output [7:0] LLKRXCHNONPOSTEDPARTIALN ;
output [7:0] LLKRXCHPOSTEDAVAILABLEN ;
output [7:0] LLKRXCHPOSTEDPARTIALN ;
output [7:0] LLKTCSTATUS ;
output [7:0] LLKTXCHCOMPLETIONREADYN ;
output [7:0] LLKTXCHNONPOSTEDREADYN ;
output [7:0] LLKTXCHPOSTEDREADYN ;
output [7:0] PIPETXDATAL0 ;
output [7:0] PIPETXDATAL1 ;
output [7:0] PIPETXDATAL2 ;
output [7:0] PIPETXDATAL3 ;
output [7:0] PIPETXDATAL4 ;
output [7:0] PIPETXDATAL5 ;
output [7:0] PIPETXDATAL6 ;
output [7:0] PIPETXDATAL7 ;
output [9:0] LLKTXCHANSPACE ;
parameter AERCAPABILITYECRCCHECKCAPABLE = "FALSE";
parameter AERCAPABILITYECRCGENCAPABLE = "FALSE";
parameter BAR0EXIST = "TRUE";
parameter BAR0PREFETCHABLE = "TRUE";
parameter BAR1EXIST = "FALSE";
parameter BAR1PREFETCHABLE = "FALSE";
parameter BAR2EXIST = "FALSE";
parameter BAR2PREFETCHABLE = "FALSE";
parameter BAR3EXIST = "FALSE";
parameter BAR3PREFETCHABLE = "FALSE";
parameter BAR4EXIST = "FALSE";
parameter BAR4PREFETCHABLE = "FALSE";
parameter BAR5EXIST = "FALSE";
parameter BAR5PREFETCHABLE = "FALSE";
parameter CLKDIVIDED = "FALSE";
parameter DUALCOREENABLE = "FALSE";
parameter DUALCORESLAVE = "FALSE";
parameter INFINITECOMPLETIONS = "TRUE";
parameter ISSWITCH = "FALSE";
parameter LINKSTATUSSLOTCLOCKCONFIG = "FALSE";
parameter LLKBYPASS = "FALSE";
parameter PBCAPABILITYSYSTEMALLOCATED = "FALSE";
parameter PCIECAPABILITYSLOTIMPL = "FALSE";
parameter PMCAPABILITYD1SUPPORT = "FALSE";
parameter PMCAPABILITYD2SUPPORT = "FALSE";
parameter PMCAPABILITYDSI = "TRUE";
parameter RAMSHARETXRX = "FALSE";
parameter RESETMODE = "FALSE";
parameter RETRYREADADDRPIPE = "FALSE";
parameter RETRYREADDATAPIPE = "FALSE";
parameter RETRYWRITEPIPE = "FALSE";
parameter RXREADADDRPIPE = "FALSE";
parameter RXREADDATAPIPE = "FALSE";
parameter RXWRITEPIPE = "FALSE";
parameter SELECTASMODE = "FALSE";
parameter SELECTDLLIF = "FALSE";
parameter SLOTCAPABILITYATTBUTTONPRESENT = "FALSE";
parameter SLOTCAPABILITYATTINDICATORPRESENT = "FALSE";
parameter SLOTCAPABILITYHOTPLUGCAPABLE = "FALSE";
parameter SLOTCAPABILITYHOTPLUGSURPRISE = "FALSE";
parameter SLOTCAPABILITYMSLSENSORPRESENT = "FALSE";
parameter SLOTCAPABILITYPOWERCONTROLLERPRESENT = "FALSE";
parameter SLOTCAPABILITYPOWERINDICATORPRESENT = "FALSE";
parameter SLOTIMPLEMENTED = "FALSE";
parameter TXREADADDRPIPE = "FALSE";
parameter TXREADDATAPIPE = "FALSE";
parameter TXWRITEPIPE = "FALSE";
parameter UPSTREAMFACING = "TRUE";
parameter XLINKSUPPORTED = "FALSE";
parameter [10:0] VC0TOTALCREDITSCD = 11'h0;
parameter [10:0] VC0TOTALCREDITSPD = 11'h34;
parameter [10:0] VC1TOTALCREDITSCD = 11'h0;
parameter [10:0] VC1TOTALCREDITSPD = 11'h0;
parameter [11:0] AERBASEPTR = 12'h110;
parameter [11:0] AERCAPABILITYNEXTPTR = 12'h138;
parameter [11:0] DSNBASEPTR = 12'h148;
parameter [11:0] DSNCAPABILITYNEXTPTR = 12'h154;
parameter [11:0] EXTCFGXPCAPPTR = 12'h0;
parameter [11:0] MSIBASEPTR = 12'h48;
parameter [11:0] PBBASEPTR = 12'h138;
parameter [11:0] PBCAPABILITYNEXTPTR = 12'h148;
parameter [11:0] PMBASEPTR = 12'h40;
parameter [11:0] RETRYRAMSIZE = 12'h9;
parameter [11:0] VCBASEPTR = 12'h154;
parameter [11:0] VCCAPABILITYNEXTPTR = 12'h0;
parameter [12:0] SLOTCAPABILITYPHYSICALSLOTNUM = 13'h0;
parameter [12:0] VC0RXFIFOBASEC = 13'h98;
parameter [12:0] VC0RXFIFOBASENP = 13'h80;
parameter [12:0] VC0RXFIFOBASEP = 13'h0;
parameter [12:0] VC0RXFIFOLIMITC = 13'h117;
parameter [12:0] VC0RXFIFOLIMITNP = 13'h97;
parameter [12:0] VC0RXFIFOLIMITP = 13'h7f;
parameter [12:0] VC0TXFIFOBASEC = 13'h98;
parameter [12:0] VC0TXFIFOBASENP = 13'h80;
parameter [12:0] VC0TXFIFOBASEP = 13'h0;
parameter [12:0] VC0TXFIFOLIMITC = 13'h117;
parameter [12:0] VC0TXFIFOLIMITNP = 13'h97;
parameter [12:0] VC0TXFIFOLIMITP = 13'h7f;
parameter [12:0] VC1RXFIFOBASEC = 13'h118;
parameter [12:0] VC1RXFIFOBASENP = 13'h118;
parameter [12:0] VC1RXFIFOBASEP = 13'h118;
parameter [12:0] VC1RXFIFOLIMITC = 13'h118;
parameter [12:0] VC1RXFIFOLIMITNP = 13'h118;
parameter [12:0] VC1RXFIFOLIMITP = 13'h118;
parameter [12:0] VC1TXFIFOBASEC = 13'h118;
parameter [12:0] VC1TXFIFOBASENP = 13'h118;
parameter [12:0] VC1TXFIFOBASEP = 13'h118;
parameter [12:0] VC1TXFIFOLIMITC = 13'h118;
parameter [12:0] VC1TXFIFOLIMITNP = 13'h118;
parameter [12:0] VC1TXFIFOLIMITP = 13'h118;
parameter [15:0] DEVICEID = 16'h5050;
parameter [15:0] SUBSYSTEMID = 16'h5050;
parameter [15:0] SUBSYSTEMVENDORID = 16'h10EE;
parameter [15:0] VENDORID = 16'h10EE;
parameter [1:0] LINKCAPABILITYASPMSUPPORT = 2'h1;
parameter [1:0] PBCAPABILITYDW0DATASCALE = 2'h0;
parameter [1:0] PBCAPABILITYDW0PMSTATE = 2'h0;
parameter [1:0] PBCAPABILITYDW1DATASCALE = 2'h0;
parameter [1:0] PBCAPABILITYDW1PMSTATE = 2'h0;
parameter [1:0] PBCAPABILITYDW2DATASCALE = 2'h0;
parameter [1:0] PBCAPABILITYDW2PMSTATE = 2'h0;
parameter [1:0] PBCAPABILITYDW3DATASCALE = 2'h0;
parameter [1:0] PBCAPABILITYDW3PMSTATE = 2'h0;
parameter [1:0] PMSTATUSCONTROLDATASCALE = 2'h0;
parameter [1:0] SLOTCAPABILITYSLOTPOWERLIMITSCALE = 2'h0;
parameter [23:0] CLASSCODE = 24'h058000;
parameter [2:0] CONFIGROUTING = 3'h1;
parameter [2:0] DEVICECAPABILITYENDPOINTL0SLATENCY = 3'h0;
parameter [2:0] DEVICECAPABILITYENDPOINTL1LATENCY = 3'h0;
parameter [2:0] MSICAPABILITYMULTIMSGCAP = 3'h0;
parameter [2:0] PBCAPABILITYDW0PMSUBSTATE = 3'h0;
parameter [2:0] PBCAPABILITYDW0POWERRAIL = 3'h0;
parameter [2:0] PBCAPABILITYDW0TYPE = 3'h0;
parameter [2:0] PBCAPABILITYDW1PMSUBSTATE = 3'h0;
parameter [2:0] PBCAPABILITYDW1POWERRAIL = 3'h0;
parameter [2:0] PBCAPABILITYDW1TYPE = 3'h0;
parameter [2:0] PBCAPABILITYDW2PMSUBSTATE = 3'h0;
parameter [2:0] PBCAPABILITYDW2POWERRAIL = 3'h0;
parameter [2:0] PBCAPABILITYDW2TYPE = 3'h0;
parameter [2:0] PBCAPABILITYDW3PMSUBSTATE = 3'h0;
parameter [2:0] PBCAPABILITYDW3POWERRAIL = 3'h0;
parameter [2:0] PBCAPABILITYDW3TYPE = 3'h0;
parameter [2:0] PMCAPABILITYAUXCURRENT = 3'h0;
parameter [2:0] PORTVCCAPABILITYEXTENDEDVCCOUNT = 3'h0;
parameter [31:0] CARDBUSCISPOINTER = 32'h0;
parameter [3:0] XPDEVICEPORTTYPE = 4'h0;
parameter [4:0] PCIECAPABILITYINTMSGNUM = 5'h0;
parameter [4:0] PMCAPABILITYPMESUPPORT = 5'h0;
parameter [5:0] BAR0MASKWIDTH = 6'h14;
parameter [5:0] BAR1MASKWIDTH = 6'h0;
parameter [5:0] BAR2MASKWIDTH = 6'h0;
parameter [5:0] BAR3MASKWIDTH = 6'h0;
parameter [5:0] BAR4MASKWIDTH = 6'h0;
parameter [5:0] BAR5MASKWIDTH = 6'h0;
parameter [5:0] LINKCAPABILITYMAXLINKWIDTH = 6'h01;
parameter [63:0] DEVICESERIALNUMBER = 64'hE000000001000A35;
parameter [6:0] VC0TOTALCREDITSCH = 7'h0;
parameter [6:0] VC0TOTALCREDITSNPH = 7'h08;
parameter [6:0] VC0TOTALCREDITSPH = 7'h08;
parameter [6:0] VC1TOTALCREDITSCH = 7'h0;
parameter [6:0] VC1TOTALCREDITSNPH = 7'h0;
parameter [6:0] VC1TOTALCREDITSPH = 7'h0;
parameter [7:0] ACTIVELANESIN = 8'h1;
parameter [7:0] CAPABILITIESPOINTER = 8'h40;
parameter [7:0] EXTCFGCAPPTR = 8'h0;
parameter [7:0] HEADERTYPE = 8'h0;
parameter [7:0] INTERRUPTPIN = 8'h0;
parameter [7:0] MSICAPABILITYNEXTPTR = 8'h60;
parameter [7:0] PBCAPABILITYDW0BASEPOWER = 8'h0;
parameter [7:0] PBCAPABILITYDW1BASEPOWER = 8'h0;
parameter [7:0] PBCAPABILITYDW2BASEPOWER = 8'h0;
parameter [7:0] PBCAPABILITYDW3BASEPOWER = 8'h0;
parameter [7:0] PCIECAPABILITYNEXTPTR = 8'h0;
parameter [7:0] PMCAPABILITYNEXTPTR = 8'h60;
parameter [7:0] PMDATA0 = 8'h0;
parameter [7:0] PMDATA1 = 8'h0;
parameter [7:0] PMDATA2 = 8'h0;
parameter [7:0] PMDATA3 = 8'h0;
parameter [7:0] PMDATA4 = 8'h0;
parameter [7:0] PMDATA5 = 8'h0;
parameter [7:0] PMDATA6 = 8'h0;
parameter [7:0] PMDATA7 = 8'h0;
parameter [7:0] PMDATA8 = 8'h0;
parameter [7:0] PORTVCCAPABILITYVCARBCAP = 8'h0;
parameter [7:0] PORTVCCAPABILITYVCARBTABLEOFFSET = 8'h0;
parameter [7:0] REVISIONID = 8'h0;
parameter [7:0] SLOTCAPABILITYSLOTPOWERLIMITVALUE = 8'h0;
parameter [7:0] XPBASEPTR = 8'h60;
parameter BAR0ADDRWIDTH = 0;
parameter BAR0IOMEMN = 0;
parameter BAR1ADDRWIDTH = 0;
parameter BAR1IOMEMN = 0;
parameter BAR2ADDRWIDTH = 0;
parameter BAR2IOMEMN = 0;
parameter BAR3ADDRWIDTH = 0;
parameter BAR3IOMEMN = 0;
parameter BAR4ADDRWIDTH = 0;
parameter BAR4IOMEMN = 0;
parameter BAR5IOMEMN = 0;
parameter DUALROLECFGCNTRLROOTEPN = 0;
parameter L0SEXITLATENCY = 7;
parameter L0SEXITLATENCYCOMCLK = 7;
parameter L1EXITLATENCY = 7;
parameter L1EXITLATENCYCOMCLK = 7;
parameter LOWPRIORITYVCCOUNT = 0;
parameter PCIEREVISION = 1;
parameter PMDATASCALE0 = 0;
parameter PMDATASCALE1 = 0;
parameter PMDATASCALE2 = 0;
parameter PMDATASCALE3 = 0;
parameter PMDATASCALE4 = 0;
parameter PMDATASCALE5 = 0;
parameter PMDATASCALE6 = 0;
parameter PMDATASCALE7 = 0;
parameter PMDATASCALE8 = 0;
parameter RETRYRAMREADLATENCY = 3;
parameter RETRYRAMWIDTH = 0;
parameter RETRYRAMWRITELATENCY = 1;
parameter TLRAMREADLATENCY = 3;
parameter TLRAMWIDTH = 0;
parameter TLRAMWRITELATENCY = 1;
parameter TXTSNFTS = 255;
parameter TXTSNFTSCOMCLK = 255;
parameter XPMAXPAYLOAD = 0;
parameter XPRCBCONTROL = 0;
endmodule
//#### END MODULE DEFINITION FOR: PCIE_INTERNAL_1_1 ####

//#### BEGIN MODULE DEFINITION FOR :PHASER_IN ###
module PHASER_IN (
  COUNTERREADVAL,
  FINEOVERFLOW,
  ICLK,
  ICLKDIV,
  ISERDESRST,
  RCLK,

  COUNTERLOADEN,
  COUNTERLOADVAL,
  COUNTERREADEN,
  DIVIDERST,
  EDGEADV,
  FINEENABLE,
  FINEINC,
  FREQREFCLK,
  MEMREFCLK,
  PHASEREFCLK,
  RANKSEL,
  RST,
  SYNCIN,
  SYSCLK
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input COUNTERLOADEN ;
input COUNTERREADEN ;
input DIVIDERST ;
input EDGEADV ;
input FINEENABLE ;
input FINEINC ;
input FREQREFCLK ;
input MEMREFCLK ;
input PHASEREFCLK ;
input RST ;
input SYNCIN ;
input SYSCLK ;
input [1:0] RANKSEL ;
input [5:0] COUNTERLOADVAL ;
output FINEOVERFLOW ;
output ICLK ;
output ICLKDIV ;
output ISERDESRST ;
output RCLK ;
output [5:0] COUNTERREADVAL ;
parameter CLKOUT_DIV = 4;
parameter DQS_BIAS_MODE = "FALSE";
parameter EN_ISERDES_RST = "FALSE";
parameter FINE_DELAY = 0;
parameter FREQ_REF_DIV = "NONE";
parameter MEMREFCLK_PERIOD = 0.000;
parameter OUTPUT_CLK_SRC = "PHASE_REF";
parameter PHASEREFCLK_PERIOD = 0.000;
parameter REFCLK_PERIOD = 0.000;
parameter SEL_CLK_OFFSET = 5;
parameter SYNC_IN_DIV_RST = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: PHASER_IN ####

//#### BEGIN MODULE DEFINITION FOR :PHASER_IN_PHY ###
module PHASER_IN_PHY (
  COUNTERREADVAL,
  DQSFOUND,
  DQSOUTOFRANGE,
  FINEOVERFLOW,
  ICLK,
  ICLKDIV,
  ISERDESRST,
  PHASELOCKED,
  RCLK,
  WRENABLE,

  BURSTPENDINGPHY,
  COUNTERLOADEN,
  COUNTERLOADVAL,
  COUNTERREADEN,
  ENCALIBPHY,
  FINEENABLE,
  FINEINC,
  FREQREFCLK,
  MEMREFCLK,
  PHASEREFCLK,
  RANKSELPHY,
  RST,
  RSTDQSFIND,
  SYNCIN,
  SYSCLK
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input BURSTPENDINGPHY ;
input COUNTERLOADEN ;
input COUNTERREADEN ;
input FINEENABLE ;
input FINEINC ;
input FREQREFCLK ;
input MEMREFCLK ;
input PHASEREFCLK ;
input RST ;
input RSTDQSFIND ;
input SYNCIN ;
input SYSCLK ;
input [1:0] ENCALIBPHY ;
input [1:0] RANKSELPHY ;
input [5:0] COUNTERLOADVAL ;
output DQSFOUND ;
output DQSOUTOFRANGE ;
output FINEOVERFLOW ;
output ICLK ;
output ICLKDIV ;
output ISERDESRST ;
output PHASELOCKED ;
output RCLK ;
output WRENABLE ;
output [5:0] COUNTERREADVAL ;
parameter BURST_MODE = "FALSE";
parameter CLKOUT_DIV = 4;
parameter [0:0] DQS_AUTO_RECAL = 1'b1;
parameter DQS_BIAS_MODE = "FALSE";
parameter [2:0] DQS_FIND_PATTERN = 3'b001;
parameter FINE_DELAY = 0;
parameter FREQ_REF_DIV = "NONE";
parameter MEMREFCLK_PERIOD = 0.000;
parameter OUTPUT_CLK_SRC = "PHASE_REF";
parameter PHASEREFCLK_PERIOD = 0.000;
parameter REFCLK_PERIOD = 0.000;
parameter SEL_CLK_OFFSET = 5;
parameter SYNC_IN_DIV_RST = "FALSE";
parameter WR_CYCLES = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: PHASER_IN_PHY ####

//#### BEGIN MODULE DEFINITION FOR :PHASER_OUT ###
module PHASER_OUT (
  COARSEOVERFLOW,
  COUNTERREADVAL,
  FINEOVERFLOW,
  OCLK,
  OCLKDELAYED,
  OCLKDIV,
  OSERDESRST,

  COARSEENABLE,
  COARSEINC,
  COUNTERLOADEN,
  COUNTERLOADVAL,
  COUNTERREADEN,
  DIVIDERST,
  EDGEADV,
  FINEENABLE,
  FINEINC,
  FREQREFCLK,
  MEMREFCLK,
  PHASEREFCLK,
  RST,
  SELFINEOCLKDELAY,
  SYNCIN,
  SYSCLK
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input COARSEENABLE ;
input COARSEINC ;
input COUNTERLOADEN ;
input COUNTERREADEN ;
input DIVIDERST ;
input EDGEADV ;
input FINEENABLE ;
input FINEINC ;
input FREQREFCLK ;
input MEMREFCLK ;
input PHASEREFCLK ;
input RST ;
input SELFINEOCLKDELAY ;
input SYNCIN ;
input SYSCLK ;
input [8:0] COUNTERLOADVAL ;
output COARSEOVERFLOW ;
output FINEOVERFLOW ;
output OCLK ;
output OCLKDELAYED ;
output OCLKDIV ;
output OSERDESRST ;
output [8:0] COUNTERREADVAL ;
parameter CLKOUT_DIV = 4;
parameter COARSE_BYPASS = "FALSE";
parameter COARSE_DELAY = 0;
parameter EN_OSERDES_RST = "FALSE";
parameter FINE_DELAY = 0;
parameter MEMREFCLK_PERIOD = 0.000;
parameter OCLKDELAY_INV = "FALSE";
parameter OCLK_DELAY = 0;
parameter OUTPUT_CLK_SRC = "PHASE_REF";
parameter PHASEREFCLK_PERIOD = 0.000;
parameter [2:0] PO = 3'b000;
parameter REFCLK_PERIOD = 0.000;
parameter SYNC_IN_DIV_RST = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: PHASER_OUT ####

//#### BEGIN MODULE DEFINITION FOR :PHASER_OUT_PHY ###
module PHASER_OUT_PHY (
  COARSEOVERFLOW,
  COUNTERREADVAL,
  CTSBUS,
  DQSBUS,
  DTSBUS,
  FINEOVERFLOW,
  OCLK,
  OCLKDELAYED,
  OCLKDIV,
  OSERDESRST,
  RDENABLE,

  BURSTPENDINGPHY,
  COARSEENABLE,
  COARSEINC,
  COUNTERLOADEN,
  COUNTERLOADVAL,
  COUNTERREADEN,
  ENCALIBPHY,
  FINEENABLE,
  FINEINC,
  FREQREFCLK,
  MEMREFCLK,
  PHASEREFCLK,
  RST,
  SELFINEOCLKDELAY,
  SYNCIN,
  SYSCLK
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input BURSTPENDINGPHY ;
input COARSEENABLE ;
input COARSEINC ;
input COUNTERLOADEN ;
input COUNTERREADEN ;
input FINEENABLE ;
input FINEINC ;
input FREQREFCLK ;
input MEMREFCLK ;
input PHASEREFCLK ;
input RST ;
input SELFINEOCLKDELAY ;
input SYNCIN ;
input SYSCLK ;
input [1:0] ENCALIBPHY ;
input [8:0] COUNTERLOADVAL ;
output COARSEOVERFLOW ;
output FINEOVERFLOW ;
output OCLK ;
output OCLKDELAYED ;
output OCLKDIV ;
output OSERDESRST ;
output RDENABLE ;
output [1:0] CTSBUS ;
output [1:0] DQSBUS ;
output [1:0] DTSBUS ;
output [8:0] COUNTERREADVAL ;
parameter CLKOUT_DIV = 4;
parameter COARSE_BYPASS = "FALSE";
parameter COARSE_DELAY = 0;
parameter DATA_CTL_N = "FALSE";
parameter DATA_RD_CYCLES = "FALSE";
parameter FINE_DELAY = 0;
parameter MEMREFCLK_PERIOD = 0.000;
parameter OCLKDELAY_INV = "FALSE";
parameter OCLK_DELAY = 0;
parameter OUTPUT_CLK_SRC = "PHASE_REF";
parameter PHASEREFCLK_PERIOD = 0.000;
parameter [2:0] PO = 3'b000;
parameter REFCLK_PERIOD = 0.000;
parameter SYNC_IN_DIV_RST = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: PHASER_OUT_PHY ####

//#### BEGIN MODULE DEFINITION FOR :PHASER_REF ###
module PHASER_REF (
  LOCKED,

  CLKIN,
  PWRDWN,
  RST
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKIN ;
input PWRDWN ;
input RST ;
output LOCKED ;
endmodule
//#### END MODULE DEFINITION FOR: PHASER_REF ####

//#### BEGIN MODULE DEFINITION FOR :PHY_CONTROL ###
module PHY_CONTROL (
  AUXOUTPUT,
  INBURSTPENDING,
  INRANKA,
  INRANKB,
  INRANKC,
  INRANKD,
  OUTBURSTPENDING,
  PCENABLECALIB,
  PHYCTLALMOSTFULL,
  PHYCTLEMPTY,
  PHYCTLFULL,
  PHYCTLREADY,

  MEMREFCLK,
  PHYCLK,
  PHYCTLMSTREMPTY,
  PHYCTLWD,
  PHYCTLWRENABLE,
  PLLLOCK,
  READCALIBENABLE,
  REFDLLLOCK,
  RESET,
  SYNCIN,
  WRITECALIBENABLE
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input MEMREFCLK ;
input PHYCLK ;
input PHYCTLMSTREMPTY ;
input PHYCTLWRENABLE ;
input PLLLOCK ;
input READCALIBENABLE ;
input REFDLLLOCK ;
input RESET ;
input SYNCIN ;
input WRITECALIBENABLE ;
input [31:0] PHYCTLWD ;
output PHYCTLALMOSTFULL ;
output PHYCTLEMPTY ;
output PHYCTLFULL ;
output PHYCTLREADY ;
output [1:0] INRANKA ;
output [1:0] INRANKB ;
output [1:0] INRANKC ;
output [1:0] INRANKD ;
output [1:0] PCENABLECALIB ;
output [3:0] AUXOUTPUT ;
output [3:0] INBURSTPENDING ;
output [3:0] OUTBURSTPENDING ;
parameter AO_TOGGLE = 0;
parameter [3:0] AO_WRLVL_EN = 4'b0000;
parameter BURST_MODE = "FALSE";
parameter CLK_RATIO = 1;
parameter CMD_OFFSET = 0;
parameter CO_DURATION = 0;
parameter DATA_CTL_A_N = "FALSE";
parameter DATA_CTL_B_N = "FALSE";
parameter DATA_CTL_C_N = "FALSE";
parameter DATA_CTL_D_N = "FALSE";
parameter DISABLE_SEQ_MATCH = "TRUE";
parameter DI_DURATION = 0;
parameter DO_DURATION = 0;
parameter EVENTS_DELAY = 63;
parameter FOUR_WINDOW_CLOCKS = 63;
parameter MULTI_REGION = "FALSE";
parameter PHY_COUNT_ENABLE = "FALSE";
parameter RD_CMD_OFFSET_0 = 0;
parameter RD_CMD_OFFSET_1 = 00;
parameter RD_CMD_OFFSET_2 = 0;
parameter RD_CMD_OFFSET_3 = 0;
parameter RD_DURATION_0 = 0;
parameter RD_DURATION_1 = 0;
parameter RD_DURATION_2 = 0;
parameter RD_DURATION_3 = 0;
parameter SYNC_MODE = "FALSE";
parameter WR_CMD_OFFSET_0 = 0;
parameter WR_CMD_OFFSET_1 = 0;
parameter WR_CMD_OFFSET_2 = 0;
parameter WR_CMD_OFFSET_3 = 0;
parameter WR_DURATION_0 = 0;
parameter WR_DURATION_1 = 0;
parameter WR_DURATION_2 = 0;
parameter WR_DURATION_3 = 0;
endmodule
//#### END MODULE DEFINITION FOR: PHY_CONTROL ####

//#### BEGIN MODULE DEFINITION FOR :PLLE2_ADV ###
module PLLE2_ADV (
  CLKFBOUT,
  CLKOUT0,
  CLKOUT1,
  CLKOUT2,
  CLKOUT3,
  CLKOUT4,
  CLKOUT5,
  DO,
  DRDY,
  LOCKED,
  CLKFBIN,
  CLKIN1,
  CLKIN2,
  CLKINSEL,
  DADDR,
  DCLK,
  DEN,
  DI,
  DWE,
  PWRDWN,
  RST
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKFBIN ;
input CLKIN1 ;
input CLKIN2 ;
input CLKINSEL ;
input DCLK ;
input DEN ;
input DWE ;
input PWRDWN ;
input RST ;
input [15:0] DI ;
input [6:0] DADDR ;
output CLKFBOUT ;
output CLKOUT0 ;
output CLKOUT1 ;
output CLKOUT2 ;
output CLKOUT3 ;
output CLKOUT4 ;
output CLKOUT5 ;
output DRDY ;
output LOCKED ;
output [15:0] DO ;
parameter BANDWIDTH = "OPTIMIZED";
parameter COMPENSATION = "ZHOLD";
parameter STARTUP_WAIT = "FALSE";
parameter CLKOUT0_DIVIDE = 1;
parameter CLKOUT1_DIVIDE = 1;
parameter CLKOUT2_DIVIDE = 1;
parameter CLKOUT3_DIVIDE = 1;
parameter CLKOUT4_DIVIDE = 1;
parameter CLKOUT5_DIVIDE = 1;
parameter DIVCLK_DIVIDE = 1;
parameter CLKFBOUT_MULT = 5;
parameter CLKFBOUT_PHASE = 0.000;
parameter CLKIN1_PERIOD = 0.000;
parameter CLKIN2_PERIOD = 0.000;
parameter CLKOUT0_DUTY_CYCLE = 0.500;
parameter CLKOUT0_PHASE = 0.000;
parameter CLKOUT1_DUTY_CYCLE = 0.500;
parameter CLKOUT1_PHASE = 0.000;
parameter CLKOUT2_DUTY_CYCLE = 0.500;
parameter CLKOUT2_PHASE = 0.000;
parameter CLKOUT3_DUTY_CYCLE = 0.500;
parameter CLKOUT3_PHASE = 0.000;
parameter CLKOUT4_DUTY_CYCLE = 0.500;
parameter CLKOUT4_PHASE = 0.000;
parameter CLKOUT5_DUTY_CYCLE = 0.500;
parameter CLKOUT5_PHASE = 0.000;
parameter REF_JITTER1 = 0.010;
parameter REF_JITTER2 = 0.010;
endmodule
//#### END MODULE DEFINITION FOR: PLLE2_ADV ####

//#### BEGIN MODULE DEFINITION FOR :PLLE2_BASE ###
module PLLE2_BASE (
  CLKFBOUT,
  CLKOUT0,
  CLKOUT1,
  CLKOUT2,
  CLKOUT3,
  CLKOUT4,
  CLKOUT5,
  LOCKED,
  CLKFBIN,
  CLKIN1,
  PWRDWN,
  RST
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKFBIN ;
input CLKIN1 ;
input PWRDWN ;
input RST ;
output CLKFBOUT ;
output CLKOUT0 ;
output CLKOUT1 ;
output CLKOUT2 ;
output CLKOUT3 ;
output CLKOUT4 ;
output CLKOUT5 ;
output LOCKED ;
parameter BANDWIDTH = "OPTIMIZED";
parameter CLKFBOUT_MULT = 5;
parameter CLKFBOUT_PHASE = 0.000;
parameter CLKIN1_PERIOD = 0.000;
parameter CLKOUT0_DIVIDE = 1;
parameter CLKOUT0_DUTY_CYCLE = 0.500;
parameter CLKOUT0_PHASE = 0.000;
parameter CLKOUT1_DIVIDE = 1;
parameter CLKOUT1_DUTY_CYCLE = 0.500;
parameter CLKOUT1_PHASE = 0.000;
parameter CLKOUT2_DIVIDE = 1;
parameter CLKOUT2_DUTY_CYCLE = 0.500;
parameter CLKOUT2_PHASE = 0.000;
parameter CLKOUT3_DIVIDE = 1;
parameter CLKOUT3_DUTY_CYCLE = 0.500;
parameter CLKOUT3_PHASE = 0.000;
parameter CLKOUT4_DIVIDE = 1;
parameter CLKOUT4_DUTY_CYCLE = 0.500;
parameter CLKOUT4_PHASE = 0.000;
parameter CLKOUT5_DIVIDE = 1;
parameter CLKOUT5_DUTY_CYCLE = 0.500;
parameter CLKOUT5_PHASE = 0.000;
parameter DIVCLK_DIVIDE = 1;
parameter REF_JITTER1 = 0.010;
parameter STARTUP_WAIT = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: PLLE2_BASE ####

//#### BEGIN MODULE DEFINITION FOR :PLL_ADV ###
module PLL_ADV (
        CLKFBDCM,
        CLKFBOUT,
        CLKOUT0,
        CLKOUT1,
        CLKOUT2,
        CLKOUT3,
        CLKOUT4,
        CLKOUT5,
        CLKOUTDCM0,
        CLKOUTDCM1,
        CLKOUTDCM2,
        CLKOUTDCM3,
        CLKOUTDCM4,
        CLKOUTDCM5,
        DO,
        DRDY,
        LOCKED,
        CLKFBIN,
        CLKIN1,
        CLKIN2,
        CLKINSEL,
        DADDR,
        DCLK,
        DEN,
        DI,
        DWE,
        REL,
        RST
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKFBIN ;
input CLKIN1 ;
input CLKIN2 ;
input CLKINSEL ;
input DCLK ;
input DEN ;
input DWE ;
input REL ;
input RST ;
input [15:0] DI ;
input [4:0] DADDR ;
output CLKFBDCM ;
output CLKFBOUT ;
output CLKOUT0 ;
output CLKOUT1 ;
output CLKOUT2 ;
output CLKOUT3 ;
output CLKOUT4 ;
output CLKOUT5 ;
output CLKOUTDCM0 ;
output CLKOUTDCM1 ;
output CLKOUTDCM2 ;
output CLKOUTDCM3 ;
output CLKOUTDCM4 ;
output CLKOUTDCM5 ;
output DRDY ;
output LOCKED ;
output [15:0] DO ;
parameter BANDWIDTH = "OPTIMIZED";
parameter CLK_FEEDBACK = "CLKFBOUT";
parameter CLKFBOUT_DESKEW_ADJUST = "NONE";
parameter CLKOUT0_DESKEW_ADJUST = "NONE";
parameter CLKOUT1_DESKEW_ADJUST = "NONE";
parameter CLKOUT2_DESKEW_ADJUST = "NONE";
parameter CLKOUT3_DESKEW_ADJUST = "NONE";
parameter CLKOUT4_DESKEW_ADJUST = "NONE";
parameter CLKOUT5_DESKEW_ADJUST = "NONE";
parameter CLKFBOUT_MULT = 1;
parameter CLKFBOUT_PHASE = 0.0;
parameter CLKIN1_PERIOD = 0.000;
parameter CLKIN2_PERIOD = 0.000;
parameter CLKOUT0_DIVIDE = 1;
parameter CLKOUT0_DUTY_CYCLE = 0.5;
parameter CLKOUT0_PHASE = 0.0;
parameter CLKOUT1_DIVIDE = 1;
parameter CLKOUT1_DUTY_CYCLE = 0.5;
parameter CLKOUT1_PHASE = 0.0;
parameter CLKOUT2_DIVIDE = 1;
parameter CLKOUT2_DUTY_CYCLE = 0.5;
parameter CLKOUT2_PHASE = 0.0;
parameter CLKOUT3_DIVIDE = 1;
parameter CLKOUT3_DUTY_CYCLE = 0.5;
parameter CLKOUT3_PHASE = 0.0;
parameter CLKOUT4_DIVIDE = 1;
parameter CLKOUT4_DUTY_CYCLE = 0.5;
parameter CLKOUT4_PHASE = 0.0;
parameter CLKOUT5_DIVIDE = 1;
parameter CLKOUT5_DUTY_CYCLE = 0.5;
parameter CLKOUT5_PHASE = 0.0;
parameter COMPENSATION = "SYSTEM_SYNCHRONOUS";
parameter DIVCLK_DIVIDE = 1;
parameter EN_REL = "FALSE";
parameter PLL_PMCD_MODE = "FALSE";
parameter REF_JITTER = 0.100;
parameter RESET_ON_LOSS_OF_LOCK = "FALSE";
parameter RST_DEASSERT_CLK = "CLKIN1";
parameter SIM_DEVICE = "VIRTEX5";
endmodule
//#### END MODULE DEFINITION FOR: PLL_ADV ####

//#### BEGIN MODULE DEFINITION FOR :PLL_BASE ###
  module PLL_BASE (
    CLKFBOUT,
    CLKOUT0,
    CLKOUT1,
    CLKOUT2,
    CLKOUT3,
    CLKOUT4,
    CLKOUT5,
    LOCKED,
    CLKFBIN,
    CLKIN,
    RST
  ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKFBIN ;
input CLKIN ;
input RST ;
output CLKFBOUT ;
output CLKOUT0 ;
output CLKOUT1 ;
output CLKOUT2 ;
output CLKOUT3 ;
output CLKOUT4 ;
output CLKOUT5 ;
output LOCKED ;
parameter BANDWIDTH = "OPTIMIZED";
parameter CLKFBOUT_MULT = 1;
parameter CLKFBOUT_PHASE = 0.0;
parameter CLKIN_PERIOD = 0.000;
parameter CLKOUT0_DIVIDE = 1;
parameter CLKOUT0_DUTY_CYCLE = 0.5;
parameter CLKOUT0_PHASE = 0.0;
parameter CLKOUT1_DIVIDE = 1;
parameter CLKOUT1_DUTY_CYCLE = 0.5;
parameter CLKOUT1_PHASE = 0.0;
parameter CLKOUT2_DIVIDE = 1;
parameter CLKOUT2_DUTY_CYCLE = 0.5;
parameter CLKOUT2_PHASE = 0.0;
parameter CLKOUT3_DIVIDE = 1;
parameter CLKOUT3_DUTY_CYCLE = 0.5;
parameter CLKOUT3_PHASE = 0.0;
parameter CLKOUT4_DIVIDE = 1;
parameter CLKOUT4_DUTY_CYCLE = 0.5;
parameter CLKOUT4_PHASE = 0.0;
parameter CLKOUT5_DIVIDE = 1;
parameter CLKOUT5_DUTY_CYCLE = 0.5;
parameter CLKOUT5_PHASE = 0.0;
parameter CLK_FEEDBACK = "CLKFBOUT";
parameter COMPENSATION = "SYSTEM_SYNCHRONOUS";
parameter DIVCLK_DIVIDE = 1;
parameter REF_JITTER = 0.100;
parameter RESET_ON_LOSS_OF_LOCK = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: PLL_BASE ####

//#### BEGIN MODULE DEFINITION FOR :PMCD ###
module PMCD (CLKA1, CLKA1D2, CLKA1D4, CLKA1D8, CLKB1, CLKC1, CLKD1, CLKA, CLKB, CLKC, CLKD, REL, RST)  /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKA ;
input CLKB ;
input CLKC ;
input CLKD ;
input REL ;
input RST ;
output CLKA1 ;
output CLKA1D2 ;
output CLKA1D4 ;
output CLKA1D8 ;
output CLKB1 ;
output CLKC1 ;
output CLKD1 ;
parameter EN_REL = "FALSE";
parameter RST_DEASSERT_CLK = "CLKA";
endmodule
//#### END MODULE DEFINITION FOR: PMCD ####

//#### BEGIN MODULE DEFINITION FOR :POST_CRC_INTERNAL ###
module POST_CRC_INTERNAL (
  CRCERROR
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
output CRCERROR ;
endmodule
//#### END MODULE DEFINITION FOR: POST_CRC_INTERNAL ####

//#### BEGIN MODULE DEFINITION FOR :PPC405_ADV ###
module PPC405_ADV (
	APUFCMDECODED,
	APUFCMDECUDI,
	APUFCMDECUDIVALID,
	APUFCMENDIAN,
	APUFCMFLUSH,
	APUFCMINSTRUCTION,
	APUFCMINSTRVALID,
	APUFCMLOADBYTEEN,
	APUFCMLOADDATA,
	APUFCMLOADDVALID,
	APUFCMOPERANDVALID,
	APUFCMRADATA,
	APUFCMRBDATA,
	APUFCMWRITEBACKOK,
	APUFCMXERCA,
	C405CPMCORESLEEPREQ,
	C405CPMMSRCE,
	C405CPMMSREE,
	C405CPMTIMERIRQ,
	C405CPMTIMERRESETREQ,
	C405DBGLOADDATAONAPUDBUS,
	C405DBGMSRWE,
	C405DBGSTOPACK,
	C405DBGWBCOMPLETE,
	C405DBGWBFULL,
	C405DBGWBIAR,
	C405JTGCAPTUREDR,
	C405JTGEXTEST,
	C405JTGPGMOUT,
	C405JTGSHIFTDR,
	C405JTGTDO,
	C405JTGTDOEN,
	C405JTGUPDATEDR,
	C405PLBDCUABORT,
	C405PLBDCUABUS,
	C405PLBDCUBE,
	C405PLBDCUCACHEABLE,
	C405PLBDCUGUARDED,
	C405PLBDCUPRIORITY,
	C405PLBDCUREQUEST,
	C405PLBDCURNW,
	C405PLBDCUSIZE2,
	C405PLBDCUU0ATTR,
	C405PLBDCUWRDBUS,
	C405PLBDCUWRITETHRU,
	C405PLBICUABORT,
	C405PLBICUABUS,
	C405PLBICUCACHEABLE,
	C405PLBICUPRIORITY,
	C405PLBICUREQUEST,
	C405PLBICUSIZE,
	C405PLBICUU0ATTR,
	C405RSTCHIPRESETREQ,
	C405RSTCORERESETREQ,
	C405RSTSYSRESETREQ,
	C405TRCCYCLE,
	C405TRCEVENEXECUTIONSTATUS,
	C405TRCODDEXECUTIONSTATUS,
	C405TRCTRACESTATUS,
	C405TRCTRIGGEREVENTOUT,
	C405TRCTRIGGEREVENTTYPE,
	C405XXXMACHINECHECK,
	DCREMACABUS,
	DCREMACCLK,
	DCREMACDBUS,
	DCREMACENABLER,
	DCREMACREAD,
	DCREMACWRITE,
	DSOCMBRAMABUS,
	DSOCMBRAMBYTEWRITE,
	DSOCMBRAMEN,
	DSOCMBRAMWRDBUS,
	DSOCMBUSY,
	DSOCMRDADDRVALID,
	DSOCMWRADDRVALID,
	EXTDCRABUS,
	EXTDCRDBUSOUT,
	EXTDCRREAD,
	EXTDCRWRITE,
	ISOCMBRAMEN,
	ISOCMBRAMEVENWRITEEN,
	ISOCMBRAMODDWRITEEN,
	ISOCMBRAMRDABUS,
	ISOCMBRAMWRABUS,
	ISOCMBRAMWRDBUS,
	ISOCMDCRBRAMEVENEN,
	ISOCMDCRBRAMODDEN,
	ISOCMDCRBRAMRDSELECT,
	BRAMDSOCMCLK,
	BRAMDSOCMRDDBUS,
	BRAMISOCMCLK,
	BRAMISOCMDCRRDDBUS,
	BRAMISOCMRDDBUS,
	CPMC405CLOCK,
	CPMC405CORECLKINACTIVE,
	CPMC405CPUCLKEN,
	CPMC405JTAGCLKEN,
	CPMC405SYNCBYPASS,
	CPMC405TIMERCLKEN,
	CPMC405TIMERTICK,
	CPMDCRCLK,
	CPMFCMCLK,
	DBGC405DEBUGHALT,
	DBGC405EXTBUSHOLDACK,
	DBGC405UNCONDDEBUGEVENT,
	DSARCVALUE,
	DSCNTLVALUE,
	DSOCMRWCOMPLETE,
	EICC405CRITINPUTIRQ,
	EICC405EXTINPUTIRQ,
	EMACDCRACK,
	EMACDCRDBUS,
	EXTDCRACK,
	EXTDCRDBUSIN,
	FCMAPUCR,
	FCMAPUDCDCREN,
	FCMAPUDCDFORCEALIGN,
	FCMAPUDCDFORCEBESTEERING,
	FCMAPUDCDFPUOP,
	FCMAPUDCDGPRWRITE,
	FCMAPUDCDLDSTBYTE,
	FCMAPUDCDLDSTDW,
	FCMAPUDCDLDSTHW,
	FCMAPUDCDLDSTQW,
	FCMAPUDCDLDSTWD,
	FCMAPUDCDLOAD,
	FCMAPUDCDPRIVOP,
	FCMAPUDCDRAEN,
	FCMAPUDCDRBEN,
	FCMAPUDCDSTORE,
	FCMAPUDCDTRAPBE,
	FCMAPUDCDTRAPLE,
	FCMAPUDCDUPDATE,
	FCMAPUDCDXERCAEN,
	FCMAPUDCDXEROVEN,
	FCMAPUDECODEBUSY,
	FCMAPUDONE,
	FCMAPUEXCEPTION,
	FCMAPUEXEBLOCKINGMCO,
	FCMAPUEXECRFIELD,
	FCMAPUEXENONBLOCKINGMCO,
	FCMAPUINSTRACK,
	FCMAPULOADWAIT,
	FCMAPURESULT,
	FCMAPURESULTVALID,
	FCMAPUSLEEPNOTREADY,
	FCMAPUXERCA,
	FCMAPUXEROV,
	ISARCVALUE,
	ISCNTLVALUE,
	JTGC405BNDSCANTDO,
	JTGC405TCK,
	JTGC405TDI,
	JTGC405TMS,
	JTGC405TRSTNEG,
	MCBCPUCLKEN,
	MCBJTAGEN,
	MCBTIMEREN,
	MCPPCRST,
	PLBC405DCUADDRACK,
	PLBC405DCUBUSY,
	PLBC405DCUERR,
	PLBC405DCURDDACK,
	PLBC405DCURDDBUS,
	PLBC405DCURDWDADDR,
	PLBC405DCUSSIZE1,
	PLBC405DCUWRDACK,
	PLBC405ICUADDRACK,
	PLBC405ICUBUSY,
	PLBC405ICUERR,
	PLBC405ICURDDACK,
	PLBC405ICURDDBUS,
	PLBC405ICURDWDADDR,
	PLBC405ICUSSIZE1,
	PLBCLK,
	RSTC405RESETCHIP,
	RSTC405RESETCORE,
	RSTC405RESETSYS,
	TIEAPUCONTROL,
	TIEAPUUDI1,
	TIEAPUUDI2,
	TIEAPUUDI3,
	TIEAPUUDI4,
	TIEAPUUDI5,
	TIEAPUUDI6,
	TIEAPUUDI7,
	TIEAPUUDI8,
	TIEC405DETERMINISTICMULT,
	TIEC405DISOPERANDFWD,
	TIEC405MMUEN,
	TIEDCRADDR,
	TIEPVRBIT10,
	TIEPVRBIT11,
	TIEPVRBIT28,
	TIEPVRBIT29,
	TIEPVRBIT30,
	TIEPVRBIT31,
	TIEPVRBIT8,
	TIEPVRBIT9,
	TRCC405TRACEDISABLE,
	TRCC405TRIGGEREVENTIN
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input BRAMDSOCMCLK ;
input BRAMISOCMCLK ;
input CPMC405CLOCK ;
input CPMC405CORECLKINACTIVE ;
input CPMC405CPUCLKEN ;
input CPMC405JTAGCLKEN ;
input CPMC405SYNCBYPASS ;
input CPMC405TIMERCLKEN ;
input CPMC405TIMERTICK ;
input CPMDCRCLK ;
input CPMFCMCLK ;
input DBGC405DEBUGHALT ;
input DBGC405EXTBUSHOLDACK ;
input DBGC405UNCONDDEBUGEVENT ;
input DSOCMRWCOMPLETE ;
input EICC405CRITINPUTIRQ ;
input EICC405EXTINPUTIRQ ;
input EMACDCRACK ;
input EXTDCRACK ;
input FCMAPUDCDCREN ;
input FCMAPUDCDFORCEALIGN ;
input FCMAPUDCDFORCEBESTEERING ;
input FCMAPUDCDFPUOP ;
input FCMAPUDCDGPRWRITE ;
input FCMAPUDCDLDSTBYTE ;
input FCMAPUDCDLDSTDW ;
input FCMAPUDCDLDSTHW ;
input FCMAPUDCDLDSTQW ;
input FCMAPUDCDLDSTWD ;
input FCMAPUDCDLOAD ;
input FCMAPUDCDPRIVOP ;
input FCMAPUDCDRAEN ;
input FCMAPUDCDRBEN ;
input FCMAPUDCDSTORE ;
input FCMAPUDCDTRAPBE ;
input FCMAPUDCDTRAPLE ;
input FCMAPUDCDUPDATE ;
input FCMAPUDCDXERCAEN ;
input FCMAPUDCDXEROVEN ;
input FCMAPUDECODEBUSY ;
input FCMAPUDONE ;
input FCMAPUEXCEPTION ;
input FCMAPUEXEBLOCKINGMCO ;
input FCMAPUEXENONBLOCKINGMCO ;
input FCMAPUINSTRACK ;
input FCMAPULOADWAIT ;
input FCMAPURESULTVALID ;
input FCMAPUSLEEPNOTREADY ;
input FCMAPUXERCA ;
input FCMAPUXEROV ;
input JTGC405BNDSCANTDO ;
input JTGC405TCK ;
input JTGC405TDI ;
input JTGC405TMS ;
input JTGC405TRSTNEG ;
input MCBCPUCLKEN ;
input MCBJTAGEN ;
input MCBTIMEREN ;
input MCPPCRST ;
input PLBC405DCUADDRACK ;
input PLBC405DCUBUSY ;
input PLBC405DCUERR ;
input PLBC405DCURDDACK ;
input PLBC405DCUSSIZE1 ;
input PLBC405DCUWRDACK ;
input PLBC405ICUADDRACK ;
input PLBC405ICUBUSY ;
input PLBC405ICUERR ;
input PLBC405ICURDDACK ;
input PLBC405ICUSSIZE1 ;
input PLBCLK ;
input RSTC405RESETCHIP ;
input RSTC405RESETCORE ;
input RSTC405RESETSYS ;
input TIEC405DETERMINISTICMULT ;
input TIEC405DISOPERANDFWD ;
input TIEC405MMUEN ;
input TIEPVRBIT10 ;
input TIEPVRBIT11 ;
input TIEPVRBIT28 ;
input TIEPVRBIT29 ;
input TIEPVRBIT30 ;
input TIEPVRBIT31 ;
input TIEPVRBIT8 ;
input TIEPVRBIT9 ;
input TRCC405TRACEDISABLE ;
input TRCC405TRIGGEREVENTIN ;
input [0:15] TIEAPUCONTROL ;
input [0:23] TIEAPUUDI1 ;
input [0:23] TIEAPUUDI2 ;
input [0:23] TIEAPUUDI3 ;
input [0:23] TIEAPUUDI4 ;
input [0:23] TIEAPUUDI5 ;
input [0:23] TIEAPUUDI6 ;
input [0:23] TIEAPUUDI7 ;
input [0:23] TIEAPUUDI8 ;
input [0:2] FCMAPUEXECRFIELD ;
input [0:31] BRAMDSOCMRDDBUS ;
input [0:31] BRAMISOCMDCRRDDBUS ;
input [0:31] EMACDCRDBUS ;
input [0:31] EXTDCRDBUSIN ;
input [0:31] FCMAPURESULT ;
input [0:3] FCMAPUCR ;
input [0:5] TIEDCRADDR ;
input [0:63] BRAMISOCMRDDBUS ;
input [0:63] PLBC405DCURDDBUS ;
input [0:63] PLBC405ICURDDBUS ;
input [0:7] DSARCVALUE ;
input [0:7] DSCNTLVALUE ;
input [0:7] ISARCVALUE ;
input [0:7] ISCNTLVALUE ;
input [1:3] PLBC405DCURDWDADDR ;
input [1:3] PLBC405ICURDWDADDR ;
output APUFCMDECODED ;
output APUFCMDECUDIVALID ;
output APUFCMENDIAN ;
output APUFCMFLUSH ;
output APUFCMINSTRVALID ;
output APUFCMLOADDVALID ;
output APUFCMOPERANDVALID ;
output APUFCMWRITEBACKOK ;
output APUFCMXERCA ;
output C405CPMCORESLEEPREQ ;
output C405CPMMSRCE ;
output C405CPMMSREE ;
output C405CPMTIMERIRQ ;
output C405CPMTIMERRESETREQ ;
output C405DBGLOADDATAONAPUDBUS ;
output C405DBGMSRWE ;
output C405DBGSTOPACK ;
output C405DBGWBCOMPLETE ;
output C405DBGWBFULL ;
output C405JTGCAPTUREDR ;
output C405JTGEXTEST ;
output C405JTGPGMOUT ;
output C405JTGSHIFTDR ;
output C405JTGTDO ;
output C405JTGTDOEN ;
output C405JTGUPDATEDR ;
output C405PLBDCUABORT ;
output C405PLBDCUCACHEABLE ;
output C405PLBDCUGUARDED ;
output C405PLBDCUREQUEST ;
output C405PLBDCURNW ;
output C405PLBDCUSIZE2 ;
output C405PLBDCUU0ATTR ;
output C405PLBDCUWRITETHRU ;
output C405PLBICUABORT ;
output C405PLBICUCACHEABLE ;
output C405PLBICUREQUEST ;
output C405PLBICUU0ATTR ;
output C405RSTCHIPRESETREQ ;
output C405RSTCORERESETREQ ;
output C405RSTSYSRESETREQ ;
output C405TRCCYCLE ;
output C405TRCTRIGGEREVENTOUT ;
output C405XXXMACHINECHECK ;
output DCREMACCLK ;
output DCREMACENABLER ;
output DCREMACREAD ;
output DCREMACWRITE ;
output DSOCMBRAMEN ;
output DSOCMBUSY ;
output DSOCMRDADDRVALID ;
output DSOCMWRADDRVALID ;
output EXTDCRREAD ;
output EXTDCRWRITE ;
output ISOCMBRAMEN ;
output ISOCMBRAMEVENWRITEEN ;
output ISOCMBRAMODDWRITEEN ;
output ISOCMDCRBRAMEVENEN ;
output ISOCMDCRBRAMODDEN ;
output ISOCMDCRBRAMRDSELECT ;
output [0:10] C405TRCTRIGGEREVENTTYPE ;
output [0:1] C405PLBDCUPRIORITY ;
output [0:1] C405PLBICUPRIORITY ;
output [0:1] C405TRCEVENEXECUTIONSTATUS ;
output [0:1] C405TRCODDEXECUTIONSTATUS ;
output [0:29] C405DBGWBIAR ;
output [0:29] C405PLBICUABUS ;
output [0:2] APUFCMDECUDI ;
output [0:31] APUFCMINSTRUCTION ;
output [0:31] APUFCMLOADDATA ;
output [0:31] APUFCMRADATA ;
output [0:31] APUFCMRBDATA ;
output [0:31] C405PLBDCUABUS ;
output [0:31] DCREMACDBUS ;
output [0:31] DSOCMBRAMWRDBUS ;
output [0:31] EXTDCRDBUSOUT ;
output [0:31] ISOCMBRAMWRDBUS ;
output [0:3] APUFCMLOADBYTEEN ;
output [0:3] C405TRCTRACESTATUS ;
output [0:3] DSOCMBRAMBYTEWRITE ;
output [0:63] C405PLBDCUWRDBUS ;
output [0:7] C405PLBDCUBE ;
output [0:9] EXTDCRABUS ;
output [2:3] C405PLBICUSIZE ;
output [8:28] ISOCMBRAMRDABUS ;
output [8:28] ISOCMBRAMWRABUS ;
output [8:29] DSOCMBRAMABUS ;
output [8:9] DCREMACABUS ;
endmodule
//#### END MODULE DEFINITION FOR: PPC405_ADV ####

//#### BEGIN MODULE DEFINITION FOR :PPC440 ###
module PPC440 (
	APUFCMDECFPUOP,
	APUFCMDECLDSTXFERSIZE,
	APUFCMDECLOAD,
	APUFCMDECNONAUTON,
	APUFCMDECSTORE,
	APUFCMDECUDI,
	APUFCMDECUDIVALID,
	APUFCMENDIAN,
	APUFCMFLUSH,
	APUFCMINSTRUCTION,
	APUFCMINSTRVALID,
	APUFCMLOADBYTEADDR,
	APUFCMLOADDATA,
	APUFCMLOADDVALID,
	APUFCMMSRFE0,
	APUFCMMSRFE1,
	APUFCMNEXTINSTRREADY,
	APUFCMOPERANDVALID,
	APUFCMRADATA,
	APUFCMRBDATA,
	APUFCMWRITEBACKOK,
	C440CPMCORESLEEPREQ,
	C440CPMDECIRPTREQ,
	C440CPMFITIRPTREQ,
	C440CPMMSRCE,
	C440CPMMSREE,
	C440CPMTIMERRESETREQ,
	C440CPMWDIRPTREQ,
	C440DBGSYSTEMCONTROL,
	C440JTGTDO,
	C440JTGTDOEN,
	C440MACHINECHECK,
	C440RSTCHIPRESETREQ,
	C440RSTCORERESETREQ,
	C440RSTSYSTEMRESETREQ,
	C440TRCBRANCHSTATUS,
	C440TRCCYCLE,
	C440TRCEXECUTIONSTATUS,
	C440TRCTRACESTATUS,
	C440TRCTRIGGEREVENTOUT,
	C440TRCTRIGGEREVENTTYPE,
	DMA0LLRSTENGINEACK,
	DMA0LLRXDSTRDYN,
	DMA0LLTXD,
	DMA0LLTXEOFN,
	DMA0LLTXEOPN,
	DMA0LLTXREM,
	DMA0LLTXSOFN,
	DMA0LLTXSOPN,
	DMA0LLTXSRCRDYN,
	DMA0RXIRQ,
	DMA0TXIRQ,
	DMA1LLRSTENGINEACK,
	DMA1LLRXDSTRDYN,
	DMA1LLTXD,
	DMA1LLTXEOFN,
	DMA1LLTXEOPN,
	DMA1LLTXREM,
	DMA1LLTXSOFN,
	DMA1LLTXSOPN,
	DMA1LLTXSRCRDYN,
	DMA1RXIRQ,
	DMA1TXIRQ,
	DMA2LLRSTENGINEACK,
	DMA2LLRXDSTRDYN,
	DMA2LLTXD,
	DMA2LLTXEOFN,
	DMA2LLTXEOPN,
	DMA2LLTXREM,
	DMA2LLTXSOFN,
	DMA2LLTXSOPN,
	DMA2LLTXSRCRDYN,
	DMA2RXIRQ,
	DMA2TXIRQ,
	DMA3LLRSTENGINEACK,
	DMA3LLRXDSTRDYN,
	DMA3LLTXD,
	DMA3LLTXEOFN,
	DMA3LLTXEOPN,
	DMA3LLTXREM,
	DMA3LLTXSOFN,
	DMA3LLTXSOPN,
	DMA3LLTXSRCRDYN,
	DMA3RXIRQ,
	DMA3TXIRQ,
	MIMCADDRESS,
	MIMCADDRESSVALID,
	MIMCBANKCONFLICT,
	MIMCBYTEENABLE,
	MIMCREADNOTWRITE,
	MIMCROWCONFLICT,
	MIMCWRITEDATA,
	MIMCWRITEDATAVALID,
	PPCCPMINTERCONNECTBUSY,
	PPCDMDCRABUS,
	PPCDMDCRDBUSOUT,
	PPCDMDCRREAD,
	PPCDMDCRUABUS,
	PPCDMDCRWRITE,
	PPCDSDCRACK,
	PPCDSDCRDBUSIN,
	PPCDSDCRTIMEOUTWAIT,
	PPCEICINTERCONNECTIRQ,
	PPCMPLBABORT,
	PPCMPLBABUS,
	PPCMPLBBE,
	PPCMPLBBUSLOCK,
	PPCMPLBLOCKERR,
	PPCMPLBPRIORITY,
	PPCMPLBRDBURST,
	PPCMPLBREQUEST,
	PPCMPLBRNW,
	PPCMPLBSIZE,
	PPCMPLBTATTRIBUTE,
	PPCMPLBTYPE,
	PPCMPLBUABUS,
	PPCMPLBWRBURST,
	PPCMPLBWRDBUS,
	PPCS0PLBADDRACK,
	PPCS0PLBMBUSY,
	PPCS0PLBMIRQ,
	PPCS0PLBMRDERR,
	PPCS0PLBMWRERR,
	PPCS0PLBRDBTERM,
	PPCS0PLBRDCOMP,
	PPCS0PLBRDDACK,
	PPCS0PLBRDDBUS,
	PPCS0PLBRDWDADDR,
	PPCS0PLBREARBITRATE,
	PPCS0PLBSSIZE,
	PPCS0PLBWAIT,
	PPCS0PLBWRBTERM,
	PPCS0PLBWRCOMP,
	PPCS0PLBWRDACK,
	PPCS1PLBADDRACK,
	PPCS1PLBMBUSY,
	PPCS1PLBMIRQ,
	PPCS1PLBMRDERR,
	PPCS1PLBMWRERR,
	PPCS1PLBRDBTERM,
	PPCS1PLBRDCOMP,
	PPCS1PLBRDDACK,
	PPCS1PLBRDDBUS,
	PPCS1PLBRDWDADDR,
	PPCS1PLBREARBITRATE,
	PPCS1PLBSSIZE,
	PPCS1PLBWAIT,
	PPCS1PLBWRBTERM,
	PPCS1PLBWRCOMP,
	PPCS1PLBWRDACK,

	CPMC440CLK,
	CPMC440CLKEN,
	CPMC440CORECLOCKINACTIVE,
	CPMC440TIMERCLOCK,
	CPMDCRCLK,
	CPMDMA0LLCLK,
	CPMDMA1LLCLK,
	CPMDMA2LLCLK,
	CPMDMA3LLCLK,
	CPMFCMCLK,
	CPMINTERCONNECTCLK,
	CPMINTERCONNECTCLKEN,
	CPMINTERCONNECTCLKNTO1,
	CPMMCCLK,
	CPMPPCMPLBCLK,
	CPMPPCS0PLBCLK,
	CPMPPCS1PLBCLK,
	DBGC440DEBUGHALT,
	DBGC440SYSTEMSTATUS,
	DBGC440UNCONDDEBUGEVENT,
	DCRPPCDMACK,
	DCRPPCDMDBUSIN,
	DCRPPCDMTIMEOUTWAIT,
	DCRPPCDSABUS,
	DCRPPCDSDBUSOUT,
	DCRPPCDSREAD,
	DCRPPCDSWRITE,
	EICC440CRITIRQ,
	EICC440EXTIRQ,
	FCMAPUCONFIRMINSTR,
	FCMAPUCR,
	FCMAPUDONE,
	FCMAPUEXCEPTION,
	FCMAPUFPSCRFEX,
	FCMAPURESULT,
	FCMAPURESULTVALID,
	FCMAPUSLEEPNOTREADY,
	FCMAPUSTOREDATA,
	JTGC440TCK,
	JTGC440TDI,
	JTGC440TMS,
	JTGC440TRSTNEG,
	LLDMA0RSTENGINEREQ,
	LLDMA0RXD,
	LLDMA0RXEOFN,
	LLDMA0RXEOPN,
	LLDMA0RXREM,
	LLDMA0RXSOFN,
	LLDMA0RXSOPN,
	LLDMA0RXSRCRDYN,
	LLDMA0TXDSTRDYN,
	LLDMA1RSTENGINEREQ,
	LLDMA1RXD,
	LLDMA1RXEOFN,
	LLDMA1RXEOPN,
	LLDMA1RXREM,
	LLDMA1RXSOFN,
	LLDMA1RXSOPN,
	LLDMA1RXSRCRDYN,
	LLDMA1TXDSTRDYN,
	LLDMA2RSTENGINEREQ,
	LLDMA2RXD,
	LLDMA2RXEOFN,
	LLDMA2RXEOPN,
	LLDMA2RXREM,
	LLDMA2RXSOFN,
	LLDMA2RXSOPN,
	LLDMA2RXSRCRDYN,
	LLDMA2TXDSTRDYN,
	LLDMA3RSTENGINEREQ,
	LLDMA3RXD,
	LLDMA3RXEOFN,
	LLDMA3RXEOPN,
	LLDMA3RXREM,
	LLDMA3RXSOFN,
	LLDMA3RXSOPN,
	LLDMA3RXSRCRDYN,
	LLDMA3TXDSTRDYN,
	MCMIADDRREADYTOACCEPT,
	MCMIREADDATA,
	MCMIREADDATAERR,
	MCMIREADDATAVALID,
	PLBPPCMADDRACK,
	PLBPPCMMBUSY,
	PLBPPCMMIRQ,
	PLBPPCMMRDERR,
	PLBPPCMMWRERR,
	PLBPPCMRDBTERM,
	PLBPPCMRDDACK,
	PLBPPCMRDDBUS,
	PLBPPCMRDPENDPRI,
	PLBPPCMRDPENDREQ,
	PLBPPCMRDWDADDR,
	PLBPPCMREARBITRATE,
	PLBPPCMREQPRI,
	PLBPPCMSSIZE,
	PLBPPCMTIMEOUT,
	PLBPPCMWRBTERM,
	PLBPPCMWRDACK,
	PLBPPCMWRPENDPRI,
	PLBPPCMWRPENDREQ,
	PLBPPCS0ABORT,
	PLBPPCS0ABUS,
	PLBPPCS0BE,
	PLBPPCS0BUSLOCK,
	PLBPPCS0LOCKERR,
	PLBPPCS0MASTERID,
	PLBPPCS0MSIZE,
	PLBPPCS0PAVALID,
	PLBPPCS0RDBURST,
	PLBPPCS0RDPENDPRI,
	PLBPPCS0RDPENDREQ,
	PLBPPCS0RDPRIM,
	PLBPPCS0REQPRI,
	PLBPPCS0RNW,
	PLBPPCS0SAVALID,
	PLBPPCS0SIZE,
	PLBPPCS0TATTRIBUTE,
	PLBPPCS0TYPE,
	PLBPPCS0UABUS,
	PLBPPCS0WRBURST,
	PLBPPCS0WRDBUS,
	PLBPPCS0WRPENDPRI,
	PLBPPCS0WRPENDREQ,
	PLBPPCS0WRPRIM,
	PLBPPCS1ABORT,
	PLBPPCS1ABUS,
	PLBPPCS1BE,
	PLBPPCS1BUSLOCK,
	PLBPPCS1LOCKERR,
	PLBPPCS1MASTERID,
	PLBPPCS1MSIZE,
	PLBPPCS1PAVALID,
	PLBPPCS1RDBURST,
	PLBPPCS1RDPENDPRI,
	PLBPPCS1RDPENDREQ,
	PLBPPCS1RDPRIM,
	PLBPPCS1REQPRI,
	PLBPPCS1RNW,
	PLBPPCS1SAVALID,
	PLBPPCS1SIZE,
	PLBPPCS1TATTRIBUTE,
	PLBPPCS1TYPE,
	PLBPPCS1UABUS,
	PLBPPCS1WRBURST,
	PLBPPCS1WRDBUS,
	PLBPPCS1WRPENDPRI,
	PLBPPCS1WRPENDREQ,
	PLBPPCS1WRPRIM,
	RSTC440RESETCHIP,
	RSTC440RESETCORE,
	RSTC440RESETSYSTEM,
	TIEC440DCURDLDCACHEPLBPRIO,
	TIEC440DCURDNONCACHEPLBPRIO,
	TIEC440DCURDTOUCHPLBPRIO,
	TIEC440DCURDURGENTPLBPRIO,
	TIEC440DCUWRFLUSHPLBPRIO,
	TIEC440DCUWRSTOREPLBPRIO,
	TIEC440DCUWRURGENTPLBPRIO,
	TIEC440ENDIANRESET,
	TIEC440ERPNRESET,
	TIEC440ICURDFETCHPLBPRIO,
	TIEC440ICURDSPECPLBPRIO,
	TIEC440ICURDTOUCHPLBPRIO,
	TIEC440PIR,
	TIEC440PVR,
	TIEC440USERRESET,
	TIEDCRBASEADDR,
	TRCC440TRACEDISABLE,
	TRCC440TRIGGEREVENTIN

) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CPMC440CLK ;
input CPMC440CLKEN ;
input CPMC440CORECLOCKINACTIVE ;
input CPMC440TIMERCLOCK ;
input CPMDCRCLK ;
input CPMDMA0LLCLK ;
input CPMDMA1LLCLK ;
input CPMDMA2LLCLK ;
input CPMDMA3LLCLK ;
input CPMFCMCLK ;
input CPMINTERCONNECTCLK ;
input CPMINTERCONNECTCLKEN ;
input CPMINTERCONNECTCLKNTO1 ;
input CPMMCCLK ;
input CPMPPCMPLBCLK ;
input CPMPPCS0PLBCLK ;
input CPMPPCS1PLBCLK ;
input DBGC440DEBUGHALT ;
input DBGC440UNCONDDEBUGEVENT ;
input DCRPPCDMACK ;
input DCRPPCDMTIMEOUTWAIT ;
input DCRPPCDSREAD ;
input DCRPPCDSWRITE ;
input EICC440CRITIRQ ;
input EICC440EXTIRQ ;
input FCMAPUCONFIRMINSTR ;
input FCMAPUDONE ;
input FCMAPUEXCEPTION ;
input FCMAPUFPSCRFEX ;
input FCMAPURESULTVALID ;
input FCMAPUSLEEPNOTREADY ;
input JTGC440TCK ;
input JTGC440TDI ;
input JTGC440TMS ;
input JTGC440TRSTNEG ;
input LLDMA0RSTENGINEREQ ;
input LLDMA0RXEOFN ;
input LLDMA0RXEOPN ;
input LLDMA0RXSOFN ;
input LLDMA0RXSOPN ;
input LLDMA0RXSRCRDYN ;
input LLDMA0TXDSTRDYN ;
input LLDMA1RSTENGINEREQ ;
input LLDMA1RXEOFN ;
input LLDMA1RXEOPN ;
input LLDMA1RXSOFN ;
input LLDMA1RXSOPN ;
input LLDMA1RXSRCRDYN ;
input LLDMA1TXDSTRDYN ;
input LLDMA2RSTENGINEREQ ;
input LLDMA2RXEOFN ;
input LLDMA2RXEOPN ;
input LLDMA2RXSOFN ;
input LLDMA2RXSOPN ;
input LLDMA2RXSRCRDYN ;
input LLDMA2TXDSTRDYN ;
input LLDMA3RSTENGINEREQ ;
input LLDMA3RXEOFN ;
input LLDMA3RXEOPN ;
input LLDMA3RXSOFN ;
input LLDMA3RXSOPN ;
input LLDMA3RXSRCRDYN ;
input LLDMA3TXDSTRDYN ;
input MCMIADDRREADYTOACCEPT ;
input MCMIREADDATAERR ;
input MCMIREADDATAVALID ;
input PLBPPCMADDRACK ;
input PLBPPCMMBUSY ;
input PLBPPCMMIRQ ;
input PLBPPCMMRDERR ;
input PLBPPCMMWRERR ;
input PLBPPCMRDBTERM ;
input PLBPPCMRDDACK ;
input PLBPPCMRDPENDREQ ;
input PLBPPCMREARBITRATE ;
input PLBPPCMTIMEOUT ;
input PLBPPCMWRBTERM ;
input PLBPPCMWRDACK ;
input PLBPPCMWRPENDREQ ;
input PLBPPCS0ABORT ;
input PLBPPCS0BUSLOCK ;
input PLBPPCS0LOCKERR ;
input PLBPPCS0PAVALID ;
input PLBPPCS0RDBURST ;
input PLBPPCS0RDPENDREQ ;
input PLBPPCS0RDPRIM ;
input PLBPPCS0RNW ;
input PLBPPCS0SAVALID ;
input PLBPPCS0WRBURST ;
input PLBPPCS0WRPENDREQ ;
input PLBPPCS0WRPRIM ;
input PLBPPCS1ABORT ;
input PLBPPCS1BUSLOCK ;
input PLBPPCS1LOCKERR ;
input PLBPPCS1PAVALID ;
input PLBPPCS1RDBURST ;
input PLBPPCS1RDPENDREQ ;
input PLBPPCS1RDPRIM ;
input PLBPPCS1RNW ;
input PLBPPCS1SAVALID ;
input PLBPPCS1WRBURST ;
input PLBPPCS1WRPENDREQ ;
input PLBPPCS1WRPRIM ;
input RSTC440RESETCHIP ;
input RSTC440RESETCORE ;
input RSTC440RESETSYSTEM ;
input TIEC440ENDIANRESET ;
input TRCC440TRACEDISABLE ;
input TRCC440TRIGGEREVENTIN ;
input [0:127] FCMAPUSTOREDATA ;
input [0:127] MCMIREADDATA ;
input [0:127] PLBPPCMRDDBUS ;
input [0:127] PLBPPCS0WRDBUS ;
input [0:127] PLBPPCS1WRDBUS ;
input [0:15] PLBPPCS0BE ;
input [0:15] PLBPPCS0TATTRIBUTE ;
input [0:15] PLBPPCS1BE ;
input [0:15] PLBPPCS1TATTRIBUTE ;
input [0:1] PLBPPCMRDPENDPRI ;
input [0:1] PLBPPCMREQPRI ;
input [0:1] PLBPPCMSSIZE ;
input [0:1] PLBPPCMWRPENDPRI ;
input [0:1] PLBPPCS0MASTERID ;
input [0:1] PLBPPCS0MSIZE ;
input [0:1] PLBPPCS0RDPENDPRI ;
input [0:1] PLBPPCS0REQPRI ;
input [0:1] PLBPPCS0WRPENDPRI ;
input [0:1] PLBPPCS1MASTERID ;
input [0:1] PLBPPCS1MSIZE ;
input [0:1] PLBPPCS1RDPENDPRI ;
input [0:1] PLBPPCS1REQPRI ;
input [0:1] PLBPPCS1WRPENDPRI ;
input [0:1] TIEC440DCURDLDCACHEPLBPRIO ;
input [0:1] TIEC440DCURDNONCACHEPLBPRIO ;
input [0:1] TIEC440DCURDTOUCHPLBPRIO ;
input [0:1] TIEC440DCURDURGENTPLBPRIO ;
input [0:1] TIEC440DCUWRFLUSHPLBPRIO ;
input [0:1] TIEC440DCUWRSTOREPLBPRIO ;
input [0:1] TIEC440DCUWRURGENTPLBPRIO ;
input [0:1] TIEC440ICURDFETCHPLBPRIO ;
input [0:1] TIEC440ICURDSPECPLBPRIO ;
input [0:1] TIEC440ICURDTOUCHPLBPRIO ;
input [0:1] TIEDCRBASEADDR ;
input [0:2] PLBPPCS0TYPE ;
input [0:2] PLBPPCS1TYPE ;
input [0:31] DCRPPCDMDBUSIN ;
input [0:31] DCRPPCDSDBUSOUT ;
input [0:31] FCMAPURESULT ;
input [0:31] LLDMA0RXD ;
input [0:31] LLDMA1RXD ;
input [0:31] LLDMA2RXD ;
input [0:31] LLDMA3RXD ;
input [0:31] PLBPPCS0ABUS ;
input [0:31] PLBPPCS1ABUS ;
input [0:3] FCMAPUCR ;
input [0:3] LLDMA0RXREM ;
input [0:3] LLDMA1RXREM ;
input [0:3] LLDMA2RXREM ;
input [0:3] LLDMA3RXREM ;
input [0:3] PLBPPCMRDWDADDR ;
input [0:3] PLBPPCS0SIZE ;
input [0:3] PLBPPCS1SIZE ;
input [0:3] TIEC440ERPNRESET ;
input [0:3] TIEC440USERRESET ;
input [0:4] DBGC440SYSTEMSTATUS ;
input [0:9] DCRPPCDSABUS ;
input [28:31] PLBPPCS0UABUS ;
input [28:31] PLBPPCS1UABUS ;
input [28:31] TIEC440PIR ;
input [28:31] TIEC440PVR ;
output APUFCMDECFPUOP ;
output APUFCMDECLOAD ;
output APUFCMDECNONAUTON ;
output APUFCMDECSTORE ;
output APUFCMDECUDIVALID ;
output APUFCMENDIAN ;
output APUFCMFLUSH ;
output APUFCMINSTRVALID ;
output APUFCMLOADDVALID ;
output APUFCMMSRFE0 ;
output APUFCMMSRFE1 ;
output APUFCMNEXTINSTRREADY ;
output APUFCMOPERANDVALID ;
output APUFCMWRITEBACKOK ;
output C440CPMCORESLEEPREQ ;
output C440CPMDECIRPTREQ ;
output C440CPMFITIRPTREQ ;
output C440CPMMSRCE ;
output C440CPMMSREE ;
output C440CPMTIMERRESETREQ ;
output C440CPMWDIRPTREQ ;
output C440JTGTDO ;
output C440JTGTDOEN ;
output C440MACHINECHECK ;
output C440RSTCHIPRESETREQ ;
output C440RSTCORERESETREQ ;
output C440RSTSYSTEMRESETREQ ;
output C440TRCCYCLE ;
output C440TRCTRIGGEREVENTOUT ;
output DMA0LLRSTENGINEACK ;
output DMA0LLRXDSTRDYN ;
output DMA0LLTXEOFN ;
output DMA0LLTXEOPN ;
output DMA0LLTXSOFN ;
output DMA0LLTXSOPN ;
output DMA0LLTXSRCRDYN ;
output DMA0RXIRQ ;
output DMA0TXIRQ ;
output DMA1LLRSTENGINEACK ;
output DMA1LLRXDSTRDYN ;
output DMA1LLTXEOFN ;
output DMA1LLTXEOPN ;
output DMA1LLTXSOFN ;
output DMA1LLTXSOPN ;
output DMA1LLTXSRCRDYN ;
output DMA1RXIRQ ;
output DMA1TXIRQ ;
output DMA2LLRSTENGINEACK ;
output DMA2LLRXDSTRDYN ;
output DMA2LLTXEOFN ;
output DMA2LLTXEOPN ;
output DMA2LLTXSOFN ;
output DMA2LLTXSOPN ;
output DMA2LLTXSRCRDYN ;
output DMA2RXIRQ ;
output DMA2TXIRQ ;
output DMA3LLRSTENGINEACK ;
output DMA3LLRXDSTRDYN ;
output DMA3LLTXEOFN ;
output DMA3LLTXEOPN ;
output DMA3LLTXSOFN ;
output DMA3LLTXSOPN ;
output DMA3LLTXSRCRDYN ;
output DMA3RXIRQ ;
output DMA3TXIRQ ;
output MIMCADDRESSVALID ;
output MIMCBANKCONFLICT ;
output MIMCREADNOTWRITE ;
output MIMCROWCONFLICT ;
output MIMCWRITEDATAVALID ;
output PPCCPMINTERCONNECTBUSY ;
output PPCDMDCRREAD ;
output PPCDMDCRWRITE ;
output PPCDSDCRACK ;
output PPCDSDCRTIMEOUTWAIT ;
output PPCEICINTERCONNECTIRQ ;
output PPCMPLBABORT ;
output PPCMPLBBUSLOCK ;
output PPCMPLBLOCKERR ;
output PPCMPLBRDBURST ;
output PPCMPLBREQUEST ;
output PPCMPLBRNW ;
output PPCMPLBWRBURST ;
output PPCS0PLBADDRACK ;
output PPCS0PLBRDBTERM ;
output PPCS0PLBRDCOMP ;
output PPCS0PLBRDDACK ;
output PPCS0PLBREARBITRATE ;
output PPCS0PLBWAIT ;
output PPCS0PLBWRBTERM ;
output PPCS0PLBWRCOMP ;
output PPCS0PLBWRDACK ;
output PPCS1PLBADDRACK ;
output PPCS1PLBRDBTERM ;
output PPCS1PLBRDCOMP ;
output PPCS1PLBRDDACK ;
output PPCS1PLBREARBITRATE ;
output PPCS1PLBWAIT ;
output PPCS1PLBWRBTERM ;
output PPCS1PLBWRCOMP ;
output PPCS1PLBWRDACK ;
output [0:127] APUFCMLOADDATA ;
output [0:127] MIMCWRITEDATA ;
output [0:127] PPCMPLBWRDBUS ;
output [0:127] PPCS0PLBRDDBUS ;
output [0:127] PPCS1PLBRDDBUS ;
output [0:13] C440TRCTRIGGEREVENTTYPE ;
output [0:15] MIMCBYTEENABLE ;
output [0:15] PPCMPLBBE ;
output [0:15] PPCMPLBTATTRIBUTE ;
output [0:1] PPCMPLBPRIORITY ;
output [0:1] PPCS0PLBSSIZE ;
output [0:1] PPCS1PLBSSIZE ;
output [0:2] APUFCMDECLDSTXFERSIZE ;
output [0:2] C440TRCBRANCHSTATUS ;
output [0:2] PPCMPLBTYPE ;
output [0:31] APUFCMINSTRUCTION ;
output [0:31] APUFCMRADATA ;
output [0:31] APUFCMRBDATA ;
output [0:31] DMA0LLTXD ;
output [0:31] DMA1LLTXD ;
output [0:31] DMA2LLTXD ;
output [0:31] DMA3LLTXD ;
output [0:31] PPCDMDCRDBUSOUT ;
output [0:31] PPCDSDCRDBUSIN ;
output [0:31] PPCMPLBABUS ;
output [0:35] MIMCADDRESS ;
output [0:3] APUFCMDECUDI ;
output [0:3] APUFCMLOADBYTEADDR ;
output [0:3] DMA0LLTXREM ;
output [0:3] DMA1LLTXREM ;
output [0:3] DMA2LLTXREM ;
output [0:3] DMA3LLTXREM ;
output [0:3] PPCMPLBSIZE ;
output [0:3] PPCS0PLBMBUSY ;
output [0:3] PPCS0PLBMIRQ ;
output [0:3] PPCS0PLBMRDERR ;
output [0:3] PPCS0PLBMWRERR ;
output [0:3] PPCS0PLBRDWDADDR ;
output [0:3] PPCS1PLBMBUSY ;
output [0:3] PPCS1PLBMIRQ ;
output [0:3] PPCS1PLBMRDERR ;
output [0:3] PPCS1PLBMWRERR ;
output [0:3] PPCS1PLBRDWDADDR ;
output [0:4] C440TRCEXECUTIONSTATUS ;
output [0:6] C440TRCTRACESTATUS ;
output [0:7] C440DBGSYSTEMCONTROL ;
output [0:9] PPCDMDCRABUS ;
output [20:21] PPCDMDCRUABUS ;
output [28:31] PPCMPLBUABUS ;
parameter CLOCK_DELAY = "FALSE";
parameter DCR_AUTOLOCK_ENABLE = "TRUE";
parameter PPCDM_ASYNCMODE = "FALSE";
parameter PPCDS_ASYNCMODE = "FALSE";
parameter PPCS0_WIDTH_128N64 = "TRUE";
parameter PPCS1_WIDTH_128N64 = "TRUE";
parameter [0:16] APU_CONTROL = 17'h02000;
parameter [0:23] APU_UDI0 = 24'h000000;
parameter [0:23] APU_UDI1 = 24'h000000;
parameter [0:23] APU_UDI10 = 24'h000000;
parameter [0:23] APU_UDI11 = 24'h000000;
parameter [0:23] APU_UDI12 = 24'h000000;
parameter [0:23] APU_UDI13 = 24'h000000;
parameter [0:23] APU_UDI14 = 24'h000000;
parameter [0:23] APU_UDI15 = 24'h000000;
parameter [0:23] APU_UDI2 = 24'h000000;
parameter [0:23] APU_UDI3 = 24'h000000;
parameter [0:23] APU_UDI4 = 24'h000000;
parameter [0:23] APU_UDI5 = 24'h000000;
parameter [0:23] APU_UDI6 = 24'h000000;
parameter [0:23] APU_UDI7 = 24'h000000;
parameter [0:23] APU_UDI8 = 24'h000000;
parameter [0:23] APU_UDI9 = 24'h000000;
parameter [0:31] DMA0_RXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA0_TXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA1_RXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA1_TXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA2_RXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA2_TXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA3_RXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA3_TXCHANNELCTRL = 32'h01010000;
parameter [0:31] INTERCONNECT_IMASK = 32'hFFFFFFFF;
parameter [0:31] INTERCONNECT_TMPL_SEL = 32'h3FFFFFFF;
parameter [0:31] MI_ARBCONFIG = 32'h00432010;
parameter [0:31] MI_BANKCONFLICT_MASK = 32'h00000000;
parameter [0:31] MI_CONTROL = 32'h0000008F;
parameter [0:31] MI_ROWCONFLICT_MASK = 32'h00000000;
parameter [0:31] PPCM_ARBCONFIG = 32'h00432010;
parameter [0:31] PPCM_CONTROL = 32'h8000009F;
parameter [0:31] PPCM_COUNTER = 32'h00000500;
parameter [0:31] PPCS0_ADDRMAP_TMPL0 = 32'hFFFFFFFF;
parameter [0:31] PPCS0_ADDRMAP_TMPL1 = 32'hFFFFFFFF;
parameter [0:31] PPCS0_ADDRMAP_TMPL2 = 32'hFFFFFFFF;
parameter [0:31] PPCS0_ADDRMAP_TMPL3 = 32'hFFFFFFFF;
parameter [0:31] PPCS0_CONTROL = 32'h8033336C;
parameter [0:31] PPCS1_ADDRMAP_TMPL0 = 32'hFFFFFFFF;
parameter [0:31] PPCS1_ADDRMAP_TMPL1 = 32'hFFFFFFFF;
parameter [0:31] PPCS1_ADDRMAP_TMPL2 = 32'hFFFFFFFF;
parameter [0:31] PPCS1_ADDRMAP_TMPL3 = 32'hFFFFFFFF;
parameter [0:31] PPCS1_CONTROL = 32'h8033336C;
parameter [0:31] XBAR_ADDRMAP_TMPL0 = 32'hFFFF0000;
parameter [0:31] XBAR_ADDRMAP_TMPL1 = 32'h00000000;
parameter [0:31] XBAR_ADDRMAP_TMPL2 = 32'h00000000;
parameter [0:31] XBAR_ADDRMAP_TMPL3 = 32'h00000000;
parameter [0:7] DMA0_CONTROL = 8'h00;
parameter [0:7] DMA1_CONTROL = 8'h00;
parameter [0:7] DMA2_CONTROL = 8'h00;
parameter [0:7] DMA3_CONTROL = 8'h00;
parameter [0:9] DMA0_RXIRQTIMER = 10'h3FF;
parameter [0:9] DMA0_TXIRQTIMER = 10'h3FF;
parameter [0:9] DMA1_RXIRQTIMER = 10'h3FF;
parameter [0:9] DMA1_TXIRQTIMER = 10'h3FF;
parameter [0:9] DMA2_RXIRQTIMER = 10'h3FF;
parameter [0:9] DMA2_TXIRQTIMER = 10'h3FF;
parameter [0:9] DMA3_RXIRQTIMER = 10'h3FF;
parameter [0:9] DMA3_TXIRQTIMER = 10'h3FF;
endmodule
//#### END MODULE DEFINITION FOR: PPC440 ####

//#### BEGIN MODULE DEFINITION FOR :PS7 ###
module PS7 (
  DMA0DATYPE,
  DMA0DAVALID,
  DMA0DRREADY,
  DMA0RSTN,
  DMA1DATYPE,
  DMA1DAVALID,
  DMA1DRREADY,
  DMA1RSTN,
  DMA2DATYPE,
  DMA2DAVALID,
  DMA2DRREADY,
  DMA2RSTN,
  DMA3DATYPE,
  DMA3DAVALID,
  DMA3DRREADY,
  DMA3RSTN,
  EMIOCAN0PHYTX,
  EMIOCAN1PHYTX,
  EMIOENET0GMIITXD,
  EMIOENET0GMIITXEN,
  EMIOENET0GMIITXER,
  EMIOENET0MDIOMDC,
  EMIOENET0MDIOO,
  EMIOENET0MDIOTN,
  EMIOENET0PTPDELAYREQRX,
  EMIOENET0PTPDELAYREQTX,
  EMIOENET0PTPPDELAYREQRX,
  EMIOENET0PTPPDELAYREQTX,
  EMIOENET0PTPPDELAYRESPRX,
  EMIOENET0PTPPDELAYRESPTX,
  EMIOENET0PTPSYNCFRAMERX,
  EMIOENET0PTPSYNCFRAMETX,
  EMIOENET0SOFRX,
  EMIOENET0SOFTX,
  EMIOENET1GMIITXD,
  EMIOENET1GMIITXEN,
  EMIOENET1GMIITXER,
  EMIOENET1MDIOMDC,
  EMIOENET1MDIOO,
  EMIOENET1MDIOTN,
  EMIOENET1PTPDELAYREQRX,
  EMIOENET1PTPDELAYREQTX,
  EMIOENET1PTPPDELAYREQRX,
  EMIOENET1PTPPDELAYREQTX,
  EMIOENET1PTPPDELAYRESPRX,
  EMIOENET1PTPPDELAYRESPTX,
  EMIOENET1PTPSYNCFRAMERX,
  EMIOENET1PTPSYNCFRAMETX,
  EMIOENET1SOFRX,
  EMIOENET1SOFTX,
  EMIOGPIOO,
  EMIOGPIOTN,
  EMIOI2C0SCLO,
  EMIOI2C0SCLTN,
  EMIOI2C0SDAO,
  EMIOI2C0SDATN,
  EMIOI2C1SCLO,
  EMIOI2C1SCLTN,
  EMIOI2C1SDAO,
  EMIOI2C1SDATN,
  EMIOPJTAGTDO,
  EMIOPJTAGTDTN,
  EMIOSDIO0BUSPOW,
  EMIOSDIO0BUSVOLT,
  EMIOSDIO0CLK,
  EMIOSDIO0CMDO,
  EMIOSDIO0CMDTN,
  EMIOSDIO0DATAO,
  EMIOSDIO0DATATN,
  EMIOSDIO0LED,
  EMIOSDIO1BUSPOW,
  EMIOSDIO1BUSVOLT,
  EMIOSDIO1CLK,
  EMIOSDIO1CMDO,
  EMIOSDIO1CMDTN,
  EMIOSDIO1DATAO,
  EMIOSDIO1DATATN,
  EMIOSDIO1LED,
  EMIOSPI0MO,
  EMIOSPI0MOTN,
  EMIOSPI0SCLKO,
  EMIOSPI0SCLKTN,
  EMIOSPI0SO,
  EMIOSPI0SSNTN,
  EMIOSPI0SSON,
  EMIOSPI0STN,
  EMIOSPI1MO,
  EMIOSPI1MOTN,
  EMIOSPI1SCLKO,
  EMIOSPI1SCLKTN,
  EMIOSPI1SO,
  EMIOSPI1SSNTN,
  EMIOSPI1SSON,
  EMIOSPI1STN,
  EMIOTRACECTL,
  EMIOTRACEDATA,
  EMIOTTC0WAVEO,
  EMIOTTC1WAVEO,
  EMIOUART0DTRN,
  EMIOUART0RTSN,
  EMIOUART0TX,
  EMIOUART1DTRN,
  EMIOUART1RTSN,
  EMIOUART1TX,
  EMIOUSB0PORTINDCTL,
  EMIOUSB0VBUSPWRSELECT,
  EMIOUSB1PORTINDCTL,
  EMIOUSB1VBUSPWRSELECT,
  EMIOWDTRSTO,
  EVENTEVENTO,
  EVENTSTANDBYWFE,
  EVENTSTANDBYWFI,
  FCLKCLK,
  FCLKRESETN,
  FTMTF2PTRIGACK,
  FTMTP2FDEBUG,
  FTMTP2FTRIG,
  IRQP2F,
  MAXIGP0ARADDR,
  MAXIGP0ARBURST,
  MAXIGP0ARCACHE,
  MAXIGP0ARESETN,
  MAXIGP0ARID,
  MAXIGP0ARLEN,
  MAXIGP0ARLOCK,
  MAXIGP0ARPROT,
  MAXIGP0ARQOS,
  MAXIGP0ARSIZE,
  MAXIGP0ARVALID,
  MAXIGP0AWADDR,
  MAXIGP0AWBURST,
  MAXIGP0AWCACHE,
  MAXIGP0AWID,
  MAXIGP0AWLEN,
  MAXIGP0AWLOCK,
  MAXIGP0AWPROT,
  MAXIGP0AWQOS,
  MAXIGP0AWSIZE,
  MAXIGP0AWVALID,
  MAXIGP0BREADY,
  MAXIGP0RREADY,
  MAXIGP0WDATA,
  MAXIGP0WID,
  MAXIGP0WLAST,
  MAXIGP0WSTRB,
  MAXIGP0WVALID,
  MAXIGP1ARADDR,
  MAXIGP1ARBURST,
  MAXIGP1ARCACHE,
  MAXIGP1ARESETN,
  MAXIGP1ARID,
  MAXIGP1ARLEN,
  MAXIGP1ARLOCK,
  MAXIGP1ARPROT,
  MAXIGP1ARQOS,
  MAXIGP1ARSIZE,
  MAXIGP1ARVALID,
  MAXIGP1AWADDR,
  MAXIGP1AWBURST,
  MAXIGP1AWCACHE,
  MAXIGP1AWID,
  MAXIGP1AWLEN,
  MAXIGP1AWLOCK,
  MAXIGP1AWPROT,
  MAXIGP1AWQOS,
  MAXIGP1AWSIZE,
  MAXIGP1AWVALID,
  MAXIGP1BREADY,
  MAXIGP1RREADY,
  MAXIGP1WDATA,
  MAXIGP1WID,
  MAXIGP1WLAST,
  MAXIGP1WSTRB,
  MAXIGP1WVALID,
  SAXIACPARESETN,
  SAXIACPARREADY,
  SAXIACPAWREADY,
  SAXIACPBID,
  SAXIACPBRESP,
  SAXIACPBVALID,
  SAXIACPRDATA,
  SAXIACPRID,
  SAXIACPRLAST,
  SAXIACPRRESP,
  SAXIACPRVALID,
  SAXIACPWREADY,
  SAXIGP0ARESETN,
  SAXIGP0ARREADY,
  SAXIGP0AWREADY,
  SAXIGP0BID,
  SAXIGP0BRESP,
  SAXIGP0BVALID,
  SAXIGP0RDATA,
  SAXIGP0RID,
  SAXIGP0RLAST,
  SAXIGP0RRESP,
  SAXIGP0RVALID,
  SAXIGP0WREADY,
  SAXIGP1ARESETN,
  SAXIGP1ARREADY,
  SAXIGP1AWREADY,
  SAXIGP1BID,
  SAXIGP1BRESP,
  SAXIGP1BVALID,
  SAXIGP1RDATA,
  SAXIGP1RID,
  SAXIGP1RLAST,
  SAXIGP1RRESP,
  SAXIGP1RVALID,
  SAXIGP1WREADY,
  SAXIHP0ARESETN,
  SAXIHP0ARREADY,
  SAXIHP0AWREADY,
  SAXIHP0BID,
  SAXIHP0BRESP,
  SAXIHP0BVALID,
  SAXIHP0RACOUNT,
  SAXIHP0RCOUNT,
  SAXIHP0RDATA,
  SAXIHP0RID,
  SAXIHP0RLAST,
  SAXIHP0RRESP,
  SAXIHP0RVALID,
  SAXIHP0WACOUNT,
  SAXIHP0WCOUNT,
  SAXIHP0WREADY,
  SAXIHP1ARESETN,
  SAXIHP1ARREADY,
  SAXIHP1AWREADY,
  SAXIHP1BID,
  SAXIHP1BRESP,
  SAXIHP1BVALID,
  SAXIHP1RACOUNT,
  SAXIHP1RCOUNT,
  SAXIHP1RDATA,
  SAXIHP1RID,
  SAXIHP1RLAST,
  SAXIHP1RRESP,
  SAXIHP1RVALID,
  SAXIHP1WACOUNT,
  SAXIHP1WCOUNT,
  SAXIHP1WREADY,
  SAXIHP2ARESETN,
  SAXIHP2ARREADY,
  SAXIHP2AWREADY,
  SAXIHP2BID,
  SAXIHP2BRESP,
  SAXIHP2BVALID,
  SAXIHP2RACOUNT,
  SAXIHP2RCOUNT,
  SAXIHP2RDATA,
  SAXIHP2RID,
  SAXIHP2RLAST,
  SAXIHP2RRESP,
  SAXIHP2RVALID,
  SAXIHP2WACOUNT,
  SAXIHP2WCOUNT,
  SAXIHP2WREADY,
  SAXIHP3ARESETN,
  SAXIHP3ARREADY,
  SAXIHP3AWREADY,
  SAXIHP3BID,
  SAXIHP3BRESP,
  SAXIHP3BVALID,
  SAXIHP3RACOUNT,
  SAXIHP3RCOUNT,
  SAXIHP3RDATA,
  SAXIHP3RID,
  SAXIHP3RLAST,
  SAXIHP3RRESP,
  SAXIHP3RVALID,
  SAXIHP3WACOUNT,
  SAXIHP3WCOUNT,
  SAXIHP3WREADY,

  DDRA,
  DDRBA,
  DDRCASB,
  DDRCKE,
  DDRCKN,
  DDRCKP,
  DDRCSB,
  DDRDM,
  DDRDQ,
  DDRDQSN,
  DDRDQSP,
  DDRDRSTB,
  DDRODT,
  DDRRASB,
  DDRVRN,
  DDRVRP,
  DDRWEB,
  MIO,
  PSCLK,
  PSPORB,
  PSSRSTB,

  DDRARB,
  DMA0ACLK,
  DMA0DAREADY,
  DMA0DRLAST,
  DMA0DRTYPE,
  DMA0DRVALID,
  DMA1ACLK,
  DMA1DAREADY,
  DMA1DRLAST,
  DMA1DRTYPE,
  DMA1DRVALID,
  DMA2ACLK,
  DMA2DAREADY,
  DMA2DRLAST,
  DMA2DRTYPE,
  DMA2DRVALID,
  DMA3ACLK,
  DMA3DAREADY,
  DMA3DRLAST,
  DMA3DRTYPE,
  DMA3DRVALID,
  EMIOCAN0PHYRX,
  EMIOCAN1PHYRX,
  EMIOENET0EXTINTIN,
  EMIOENET0GMIICOL,
  EMIOENET0GMIICRS,
  EMIOENET0GMIIRXCLK,
  EMIOENET0GMIIRXD,
  EMIOENET0GMIIRXDV,
  EMIOENET0GMIIRXER,
  EMIOENET0GMIITXCLK,
  EMIOENET0MDIOI,
  EMIOENET1EXTINTIN,
  EMIOENET1GMIICOL,
  EMIOENET1GMIICRS,
  EMIOENET1GMIIRXCLK,
  EMIOENET1GMIIRXD,
  EMIOENET1GMIIRXDV,
  EMIOENET1GMIIRXER,
  EMIOENET1GMIITXCLK,
  EMIOENET1MDIOI,
  EMIOGPIOI,
  EMIOI2C0SCLI,
  EMIOI2C0SDAI,
  EMIOI2C1SCLI,
  EMIOI2C1SDAI,
  EMIOPJTAGTCK,
  EMIOPJTAGTDI,
  EMIOPJTAGTMS,
  EMIOSDIO0CDN,
  EMIOSDIO0CLKFB,
  EMIOSDIO0CMDI,
  EMIOSDIO0DATAI,
  EMIOSDIO0WP,
  EMIOSDIO1CDN,
  EMIOSDIO1CLKFB,
  EMIOSDIO1CMDI,
  EMIOSDIO1DATAI,
  EMIOSDIO1WP,
  EMIOSPI0MI,
  EMIOSPI0SCLKI,
  EMIOSPI0SI,
  EMIOSPI0SSIN,
  EMIOSPI1MI,
  EMIOSPI1SCLKI,
  EMIOSPI1SI,
  EMIOSPI1SSIN,
  EMIOSRAMINTIN,
  EMIOTRACECLK,
  EMIOTTC0CLKI,
  EMIOTTC1CLKI,
  EMIOUART0CTSN,
  EMIOUART0DCDN,
  EMIOUART0DSRN,
  EMIOUART0RIN,
  EMIOUART0RX,
  EMIOUART1CTSN,
  EMIOUART1DCDN,
  EMIOUART1DSRN,
  EMIOUART1RIN,
  EMIOUART1RX,
  EMIOUSB0VBUSPWRFAULT,
  EMIOUSB1VBUSPWRFAULT,
  EMIOWDTCLKI,
  EVENTEVENTI,
  FCLKCLKTRIGN,
  FPGAIDLEN,
  FTMDTRACEINATID,
  FTMDTRACEINCLOCK,
  FTMDTRACEINDATA,
  FTMDTRACEINVALID,
  FTMTF2PDEBUG,
  FTMTF2PTRIG,
  FTMTP2FTRIGACK,
  IRQF2P,
  MAXIGP0ACLK,
  MAXIGP0ARREADY,
  MAXIGP0AWREADY,
  MAXIGP0BID,
  MAXIGP0BRESP,
  MAXIGP0BVALID,
  MAXIGP0RDATA,
  MAXIGP0RID,
  MAXIGP0RLAST,
  MAXIGP0RRESP,
  MAXIGP0RVALID,
  MAXIGP0WREADY,
  MAXIGP1ACLK,
  MAXIGP1ARREADY,
  MAXIGP1AWREADY,
  MAXIGP1BID,
  MAXIGP1BRESP,
  MAXIGP1BVALID,
  MAXIGP1RDATA,
  MAXIGP1RID,
  MAXIGP1RLAST,
  MAXIGP1RRESP,
  MAXIGP1RVALID,
  MAXIGP1WREADY,
  SAXIACPACLK,
  SAXIACPARADDR,
  SAXIACPARBURST,
  SAXIACPARCACHE,
  SAXIACPARID,
  SAXIACPARLEN,
  SAXIACPARLOCK,
  SAXIACPARPROT,
  SAXIACPARQOS,
  SAXIACPARSIZE,
  SAXIACPARUSER,
  SAXIACPARVALID,
  SAXIACPAWADDR,
  SAXIACPAWBURST,
  SAXIACPAWCACHE,
  SAXIACPAWID,
  SAXIACPAWLEN,
  SAXIACPAWLOCK,
  SAXIACPAWPROT,
  SAXIACPAWQOS,
  SAXIACPAWSIZE,
  SAXIACPAWUSER,
  SAXIACPAWVALID,
  SAXIACPBREADY,
  SAXIACPRREADY,
  SAXIACPWDATA,
  SAXIACPWID,
  SAXIACPWLAST,
  SAXIACPWSTRB,
  SAXIACPWVALID,
  SAXIGP0ACLK,
  SAXIGP0ARADDR,
  SAXIGP0ARBURST,
  SAXIGP0ARCACHE,
  SAXIGP0ARID,
  SAXIGP0ARLEN,
  SAXIGP0ARLOCK,
  SAXIGP0ARPROT,
  SAXIGP0ARQOS,
  SAXIGP0ARSIZE,
  SAXIGP0ARVALID,
  SAXIGP0AWADDR,
  SAXIGP0AWBURST,
  SAXIGP0AWCACHE,
  SAXIGP0AWID,
  SAXIGP0AWLEN,
  SAXIGP0AWLOCK,
  SAXIGP0AWPROT,
  SAXIGP0AWQOS,
  SAXIGP0AWSIZE,
  SAXIGP0AWVALID,
  SAXIGP0BREADY,
  SAXIGP0RREADY,
  SAXIGP0WDATA,
  SAXIGP0WID,
  SAXIGP0WLAST,
  SAXIGP0WSTRB,
  SAXIGP0WVALID,
  SAXIGP1ACLK,
  SAXIGP1ARADDR,
  SAXIGP1ARBURST,
  SAXIGP1ARCACHE,
  SAXIGP1ARID,
  SAXIGP1ARLEN,
  SAXIGP1ARLOCK,
  SAXIGP1ARPROT,
  SAXIGP1ARQOS,
  SAXIGP1ARSIZE,
  SAXIGP1ARVALID,
  SAXIGP1AWADDR,
  SAXIGP1AWBURST,
  SAXIGP1AWCACHE,
  SAXIGP1AWID,
  SAXIGP1AWLEN,
  SAXIGP1AWLOCK,
  SAXIGP1AWPROT,
  SAXIGP1AWQOS,
  SAXIGP1AWSIZE,
  SAXIGP1AWVALID,
  SAXIGP1BREADY,
  SAXIGP1RREADY,
  SAXIGP1WDATA,
  SAXIGP1WID,
  SAXIGP1WLAST,
  SAXIGP1WSTRB,
  SAXIGP1WVALID,
  SAXIHP0ACLK,
  SAXIHP0ARADDR,
  SAXIHP0ARBURST,
  SAXIHP0ARCACHE,
  SAXIHP0ARID,
  SAXIHP0ARLEN,
  SAXIHP0ARLOCK,
  SAXIHP0ARPROT,
  SAXIHP0ARQOS,
  SAXIHP0ARSIZE,
  SAXIHP0ARVALID,
  SAXIHP0AWADDR,
  SAXIHP0AWBURST,
  SAXIHP0AWCACHE,
  SAXIHP0AWID,
  SAXIHP0AWLEN,
  SAXIHP0AWLOCK,
  SAXIHP0AWPROT,
  SAXIHP0AWQOS,
  SAXIHP0AWSIZE,
  SAXIHP0AWVALID,
  SAXIHP0BREADY,
  SAXIHP0RDISSUECAP1EN,
  SAXIHP0RREADY,
  SAXIHP0WDATA,
  SAXIHP0WID,
  SAXIHP0WLAST,
  SAXIHP0WRISSUECAP1EN,
  SAXIHP0WSTRB,
  SAXIHP0WVALID,
  SAXIHP1ACLK,
  SAXIHP1ARADDR,
  SAXIHP1ARBURST,
  SAXIHP1ARCACHE,
  SAXIHP1ARID,
  SAXIHP1ARLEN,
  SAXIHP1ARLOCK,
  SAXIHP1ARPROT,
  SAXIHP1ARQOS,
  SAXIHP1ARSIZE,
  SAXIHP1ARVALID,
  SAXIHP1AWADDR,
  SAXIHP1AWBURST,
  SAXIHP1AWCACHE,
  SAXIHP1AWID,
  SAXIHP1AWLEN,
  SAXIHP1AWLOCK,
  SAXIHP1AWPROT,
  SAXIHP1AWQOS,
  SAXIHP1AWSIZE,
  SAXIHP1AWVALID,
  SAXIHP1BREADY,
  SAXIHP1RDISSUECAP1EN,
  SAXIHP1RREADY,
  SAXIHP1WDATA,
  SAXIHP1WID,
  SAXIHP1WLAST,
  SAXIHP1WRISSUECAP1EN,
  SAXIHP1WSTRB,
  SAXIHP1WVALID,
  SAXIHP2ACLK,
  SAXIHP2ARADDR,
  SAXIHP2ARBURST,
  SAXIHP2ARCACHE,
  SAXIHP2ARID,
  SAXIHP2ARLEN,
  SAXIHP2ARLOCK,
  SAXIHP2ARPROT,
  SAXIHP2ARQOS,
  SAXIHP2ARSIZE,
  SAXIHP2ARVALID,
  SAXIHP2AWADDR,
  SAXIHP2AWBURST,
  SAXIHP2AWCACHE,
  SAXIHP2AWID,
  SAXIHP2AWLEN,
  SAXIHP2AWLOCK,
  SAXIHP2AWPROT,
  SAXIHP2AWQOS,
  SAXIHP2AWSIZE,
  SAXIHP2AWVALID,
  SAXIHP2BREADY,
  SAXIHP2RDISSUECAP1EN,
  SAXIHP2RREADY,
  SAXIHP2WDATA,
  SAXIHP2WID,
  SAXIHP2WLAST,
  SAXIHP2WRISSUECAP1EN,
  SAXIHP2WSTRB,
  SAXIHP2WVALID,
  SAXIHP3ACLK,
  SAXIHP3ARADDR,
  SAXIHP3ARBURST,
  SAXIHP3ARCACHE,
  SAXIHP3ARID,
  SAXIHP3ARLEN,
  SAXIHP3ARLOCK,
  SAXIHP3ARPROT,
  SAXIHP3ARQOS,
  SAXIHP3ARSIZE,
  SAXIHP3ARVALID,
  SAXIHP3AWADDR,
  SAXIHP3AWBURST,
  SAXIHP3AWCACHE,
  SAXIHP3AWID,
  SAXIHP3AWLEN,
  SAXIHP3AWLOCK,
  SAXIHP3AWPROT,
  SAXIHP3AWQOS,
  SAXIHP3AWSIZE,
  SAXIHP3AWVALID,
  SAXIHP3BREADY,
  SAXIHP3RDISSUECAP1EN,
  SAXIHP3RREADY,
  SAXIHP3WDATA,
  SAXIHP3WID,
  SAXIHP3WLAST,
  SAXIHP3WRISSUECAP1EN,
  SAXIHP3WSTRB,
  SAXIHP3WVALID
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input DMA0ACLK ;
input DMA0DAREADY ;
input DMA0DRLAST ;
input DMA0DRVALID ;
input DMA1ACLK ;
input DMA1DAREADY ;
input DMA1DRLAST ;
input DMA1DRVALID ;
input DMA2ACLK ;
input DMA2DAREADY ;
input DMA2DRLAST ;
input DMA2DRVALID ;
input DMA3ACLK ;
input DMA3DAREADY ;
input DMA3DRLAST ;
input DMA3DRVALID ;
input EMIOCAN0PHYRX ;
input EMIOCAN1PHYRX ;
input EMIOENET0EXTINTIN ;
input EMIOENET0GMIICOL ;
input EMIOENET0GMIICRS ;
input EMIOENET0GMIIRXCLK ;
input EMIOENET0GMIIRXDV ;
input EMIOENET0GMIIRXER ;
input EMIOENET0GMIITXCLK ;
input EMIOENET0MDIOI ;
input EMIOENET1EXTINTIN ;
input EMIOENET1GMIICOL ;
input EMIOENET1GMIICRS ;
input EMIOENET1GMIIRXCLK ;
input EMIOENET1GMIIRXDV ;
input EMIOENET1GMIIRXER ;
input EMIOENET1GMIITXCLK ;
input EMIOENET1MDIOI ;
input EMIOI2C0SCLI ;
input EMIOI2C0SDAI ;
input EMIOI2C1SCLI ;
input EMIOI2C1SDAI ;
input EMIOPJTAGTCK ;
input EMIOPJTAGTDI ;
input EMIOPJTAGTMS ;
input EMIOSDIO0CDN ;
input EMIOSDIO0CLKFB ;
input EMIOSDIO0CMDI ;
input EMIOSDIO0WP ;
input EMIOSDIO1CDN ;
input EMIOSDIO1CLKFB ;
input EMIOSDIO1CMDI ;
input EMIOSDIO1WP ;
input EMIOSPI0MI ;
input EMIOSPI0SCLKI ;
input EMIOSPI0SI ;
input EMIOSPI0SSIN ;
input EMIOSPI1MI ;
input EMIOSPI1SCLKI ;
input EMIOSPI1SI ;
input EMIOSPI1SSIN ;
input EMIOSRAMINTIN ;
input EMIOTRACECLK ;
input EMIOUART0CTSN ;
input EMIOUART0DCDN ;
input EMIOUART0DSRN ;
input EMIOUART0RIN ;
input EMIOUART0RX ;
input EMIOUART1CTSN ;
input EMIOUART1DCDN ;
input EMIOUART1DSRN ;
input EMIOUART1RIN ;
input EMIOUART1RX ;
input EMIOUSB0VBUSPWRFAULT ;
input EMIOUSB1VBUSPWRFAULT ;
input EMIOWDTCLKI ;
input EVENTEVENTI ;
input FPGAIDLEN ;
input FTMDTRACEINCLOCK ;
input FTMDTRACEINVALID ;
input MAXIGP0ACLK ;
input MAXIGP0ARREADY ;
input MAXIGP0AWREADY ;
input MAXIGP0BVALID ;
input MAXIGP0RLAST ;
input MAXIGP0RVALID ;
input MAXIGP0WREADY ;
input MAXIGP1ACLK ;
input MAXIGP1ARREADY ;
input MAXIGP1AWREADY ;
input MAXIGP1BVALID ;
input MAXIGP1RLAST ;
input MAXIGP1RVALID ;
input MAXIGP1WREADY ;
input SAXIACPACLK ;
input SAXIACPARVALID ;
input SAXIACPAWVALID ;
input SAXIACPBREADY ;
input SAXIACPRREADY ;
input SAXIACPWLAST ;
input SAXIACPWVALID ;
input SAXIGP0ACLK ;
input SAXIGP0ARVALID ;
input SAXIGP0AWVALID ;
input SAXIGP0BREADY ;
input SAXIGP0RREADY ;
input SAXIGP0WLAST ;
input SAXIGP0WVALID ;
input SAXIGP1ACLK ;
input SAXIGP1ARVALID ;
input SAXIGP1AWVALID ;
input SAXIGP1BREADY ;
input SAXIGP1RREADY ;
input SAXIGP1WLAST ;
input SAXIGP1WVALID ;
input SAXIHP0ACLK ;
input SAXIHP0ARVALID ;
input SAXIHP0AWVALID ;
input SAXIHP0BREADY ;
input SAXIHP0RDISSUECAP1EN ;
input SAXIHP0RREADY ;
input SAXIHP0WLAST ;
input SAXIHP0WRISSUECAP1EN ;
input SAXIHP0WVALID ;
input SAXIHP1ACLK ;
input SAXIHP1ARVALID ;
input SAXIHP1AWVALID ;
input SAXIHP1BREADY ;
input SAXIHP1RDISSUECAP1EN ;
input SAXIHP1RREADY ;
input SAXIHP1WLAST ;
input SAXIHP1WRISSUECAP1EN ;
input SAXIHP1WVALID ;
input SAXIHP2ACLK ;
input SAXIHP2ARVALID ;
input SAXIHP2AWVALID ;
input SAXIHP2BREADY ;
input SAXIHP2RDISSUECAP1EN ;
input SAXIHP2RREADY ;
input SAXIHP2WLAST ;
input SAXIHP2WRISSUECAP1EN ;
input SAXIHP2WVALID ;
input SAXIHP3ACLK ;
input SAXIHP3ARVALID ;
input SAXIHP3AWVALID ;
input SAXIHP3BREADY ;
input SAXIHP3RDISSUECAP1EN ;
input SAXIHP3RREADY ;
input SAXIHP3WLAST ;
input SAXIHP3WRISSUECAP1EN ;
input SAXIHP3WVALID ;
input [11:0] MAXIGP0BID ;
input [11:0] MAXIGP0RID ;
input [11:0] MAXIGP1BID ;
input [11:0] MAXIGP1RID ;
input [19:0] IRQF2P ;
input [1:0] DMA0DRTYPE ;
input [1:0] DMA1DRTYPE ;
input [1:0] DMA2DRTYPE ;
input [1:0] DMA3DRTYPE ;
input [1:0] MAXIGP0BRESP ;
input [1:0] MAXIGP0RRESP ;
input [1:0] MAXIGP1BRESP ;
input [1:0] MAXIGP1RRESP ;
input [1:0] SAXIACPARBURST ;
input [1:0] SAXIACPARLOCK ;
input [1:0] SAXIACPARSIZE ;
input [1:0] SAXIACPAWBURST ;
input [1:0] SAXIACPAWLOCK ;
input [1:0] SAXIACPAWSIZE ;
input [1:0] SAXIGP0ARBURST ;
input [1:0] SAXIGP0ARLOCK ;
input [1:0] SAXIGP0ARSIZE ;
input [1:0] SAXIGP0AWBURST ;
input [1:0] SAXIGP0AWLOCK ;
input [1:0] SAXIGP0AWSIZE ;
input [1:0] SAXIGP1ARBURST ;
input [1:0] SAXIGP1ARLOCK ;
input [1:0] SAXIGP1ARSIZE ;
input [1:0] SAXIGP1AWBURST ;
input [1:0] SAXIGP1AWLOCK ;
input [1:0] SAXIGP1AWSIZE ;
input [1:0] SAXIHP0ARBURST ;
input [1:0] SAXIHP0ARLOCK ;
input [1:0] SAXIHP0ARSIZE ;
input [1:0] SAXIHP0AWBURST ;
input [1:0] SAXIHP0AWLOCK ;
input [1:0] SAXIHP0AWSIZE ;
input [1:0] SAXIHP1ARBURST ;
input [1:0] SAXIHP1ARLOCK ;
input [1:0] SAXIHP1ARSIZE ;
input [1:0] SAXIHP1AWBURST ;
input [1:0] SAXIHP1AWLOCK ;
input [1:0] SAXIHP1AWSIZE ;
input [1:0] SAXIHP2ARBURST ;
input [1:0] SAXIHP2ARLOCK ;
input [1:0] SAXIHP2ARSIZE ;
input [1:0] SAXIHP2AWBURST ;
input [1:0] SAXIHP2AWLOCK ;
input [1:0] SAXIHP2AWSIZE ;
input [1:0] SAXIHP3ARBURST ;
input [1:0] SAXIHP3ARLOCK ;
input [1:0] SAXIHP3ARSIZE ;
input [1:0] SAXIHP3AWBURST ;
input [1:0] SAXIHP3AWLOCK ;
input [1:0] SAXIHP3AWSIZE ;
input [2:0] EMIOTTC0CLKI ;
input [2:0] EMIOTTC1CLKI ;
input [2:0] SAXIACPARID ;
input [2:0] SAXIACPARPROT ;
input [2:0] SAXIACPAWID ;
input [2:0] SAXIACPAWPROT ;
input [2:0] SAXIACPWID ;
input [2:0] SAXIGP0ARPROT ;
input [2:0] SAXIGP0AWPROT ;
input [2:0] SAXIGP1ARPROT ;
input [2:0] SAXIGP1AWPROT ;
input [2:0] SAXIHP0ARPROT ;
input [2:0] SAXIHP0AWPROT ;
input [2:0] SAXIHP1ARPROT ;
input [2:0] SAXIHP1AWPROT ;
input [2:0] SAXIHP2ARPROT ;
input [2:0] SAXIHP2AWPROT ;
input [2:0] SAXIHP3ARPROT ;
input [2:0] SAXIHP3AWPROT ;
input [31:0] FTMDTRACEINDATA ;
input [31:0] FTMTF2PDEBUG ;
input [31:0] MAXIGP0RDATA ;
input [31:0] MAXIGP1RDATA ;
input [31:0] SAXIACPARADDR ;
input [31:0] SAXIACPAWADDR ;
input [31:0] SAXIGP0ARADDR ;
input [31:0] SAXIGP0AWADDR ;
input [31:0] SAXIGP0WDATA ;
input [31:0] SAXIGP1ARADDR ;
input [31:0] SAXIGP1AWADDR ;
input [31:0] SAXIGP1WDATA ;
input [31:0] SAXIHP0ARADDR ;
input [31:0] SAXIHP0AWADDR ;
input [31:0] SAXIHP1ARADDR ;
input [31:0] SAXIHP1AWADDR ;
input [31:0] SAXIHP2ARADDR ;
input [31:0] SAXIHP2AWADDR ;
input [31:0] SAXIHP3ARADDR ;
input [31:0] SAXIHP3AWADDR ;
input [3:0] DDRARB ;
input [3:0] EMIOSDIO0DATAI ;
input [3:0] EMIOSDIO1DATAI ;
input [3:0] FCLKCLKTRIGN ;
input [3:0] FTMDTRACEINATID ;
input [3:0] FTMTF2PTRIG ;
input [3:0] FTMTP2FTRIGACK ;
input [3:0] SAXIACPARCACHE ;
input [3:0] SAXIACPARLEN ;
input [3:0] SAXIACPARQOS ;
input [3:0] SAXIACPAWCACHE ;
input [3:0] SAXIACPAWLEN ;
input [3:0] SAXIACPAWQOS ;
input [3:0] SAXIGP0ARCACHE ;
input [3:0] SAXIGP0ARLEN ;
input [3:0] SAXIGP0ARQOS ;
input [3:0] SAXIGP0AWCACHE ;
input [3:0] SAXIGP0AWLEN ;
input [3:0] SAXIGP0AWQOS ;
input [3:0] SAXIGP0WSTRB ;
input [3:0] SAXIGP1ARCACHE ;
input [3:0] SAXIGP1ARLEN ;
input [3:0] SAXIGP1ARQOS ;
input [3:0] SAXIGP1AWCACHE ;
input [3:0] SAXIGP1AWLEN ;
input [3:0] SAXIGP1AWQOS ;
input [3:0] SAXIGP1WSTRB ;
input [3:0] SAXIHP0ARCACHE ;
input [3:0] SAXIHP0ARLEN ;
input [3:0] SAXIHP0ARQOS ;
input [3:0] SAXIHP0AWCACHE ;
input [3:0] SAXIHP0AWLEN ;
input [3:0] SAXIHP0AWQOS ;
input [3:0] SAXIHP1ARCACHE ;
input [3:0] SAXIHP1ARLEN ;
input [3:0] SAXIHP1ARQOS ;
input [3:0] SAXIHP1AWCACHE ;
input [3:0] SAXIHP1AWLEN ;
input [3:0] SAXIHP1AWQOS ;
input [3:0] SAXIHP2ARCACHE ;
input [3:0] SAXIHP2ARLEN ;
input [3:0] SAXIHP2ARQOS ;
input [3:0] SAXIHP2AWCACHE ;
input [3:0] SAXIHP2AWLEN ;
input [3:0] SAXIHP2AWQOS ;
input [3:0] SAXIHP3ARCACHE ;
input [3:0] SAXIHP3ARLEN ;
input [3:0] SAXIHP3ARQOS ;
input [3:0] SAXIHP3AWCACHE ;
input [3:0] SAXIHP3AWLEN ;
input [3:0] SAXIHP3AWQOS ;
input [4:0] SAXIACPARUSER ;
input [4:0] SAXIACPAWUSER ;
input [5:0] SAXIGP0ARID ;
input [5:0] SAXIGP0AWID ;
input [5:0] SAXIGP0WID ;
input [5:0] SAXIGP1ARID ;
input [5:0] SAXIGP1AWID ;
input [5:0] SAXIGP1WID ;
input [5:0] SAXIHP0ARID ;
input [5:0] SAXIHP0AWID ;
input [5:0] SAXIHP0WID ;
input [5:0] SAXIHP1ARID ;
input [5:0] SAXIHP1AWID ;
input [5:0] SAXIHP1WID ;
input [5:0] SAXIHP2ARID ;
input [5:0] SAXIHP2AWID ;
input [5:0] SAXIHP2WID ;
input [5:0] SAXIHP3ARID ;
input [5:0] SAXIHP3AWID ;
input [5:0] SAXIHP3WID ;
input [63:0] EMIOGPIOI ;
input [63:0] SAXIACPWDATA ;
input [63:0] SAXIHP0WDATA ;
input [63:0] SAXIHP1WDATA ;
input [63:0] SAXIHP2WDATA ;
input [63:0] SAXIHP3WDATA ;
input [7:0] EMIOENET0GMIIRXD ;
input [7:0] EMIOENET1GMIIRXD ;
input [7:0] SAXIACPWSTRB ;
input [7:0] SAXIHP0WSTRB ;
input [7:0] SAXIHP1WSTRB ;
input [7:0] SAXIHP2WSTRB ;
input [7:0] SAXIHP3WSTRB ;
output DMA0DAVALID ;
output DMA0DRREADY ;
output DMA0RSTN ;
output DMA1DAVALID ;
output DMA1DRREADY ;
output DMA1RSTN ;
output DMA2DAVALID ;
output DMA2DRREADY ;
output DMA2RSTN ;
output DMA3DAVALID ;
output DMA3DRREADY ;
output DMA3RSTN ;
output EMIOCAN0PHYTX ;
output EMIOCAN1PHYTX ;
output EMIOENET0GMIITXEN ;
output EMIOENET0GMIITXER ;
output EMIOENET0MDIOMDC ;
output EMIOENET0MDIOO ;
output EMIOENET0MDIOTN ;
output EMIOENET0PTPDELAYREQRX ;
output EMIOENET0PTPDELAYREQTX ;
output EMIOENET0PTPPDELAYREQRX ;
output EMIOENET0PTPPDELAYREQTX ;
output EMIOENET0PTPPDELAYRESPRX ;
output EMIOENET0PTPPDELAYRESPTX ;
output EMIOENET0PTPSYNCFRAMERX ;
output EMIOENET0PTPSYNCFRAMETX ;
output EMIOENET0SOFRX ;
output EMIOENET0SOFTX ;
output EMIOENET1GMIITXEN ;
output EMIOENET1GMIITXER ;
output EMIOENET1MDIOMDC ;
output EMIOENET1MDIOO ;
output EMIOENET1MDIOTN ;
output EMIOENET1PTPDELAYREQRX ;
output EMIOENET1PTPDELAYREQTX ;
output EMIOENET1PTPPDELAYREQRX ;
output EMIOENET1PTPPDELAYREQTX ;
output EMIOENET1PTPPDELAYRESPRX ;
output EMIOENET1PTPPDELAYRESPTX ;
output EMIOENET1PTPSYNCFRAMERX ;
output EMIOENET1PTPSYNCFRAMETX ;
output EMIOENET1SOFRX ;
output EMIOENET1SOFTX ;
output EMIOI2C0SCLO ;
output EMIOI2C0SCLTN ;
output EMIOI2C0SDAO ;
output EMIOI2C0SDATN ;
output EMIOI2C1SCLO ;
output EMIOI2C1SCLTN ;
output EMIOI2C1SDAO ;
output EMIOI2C1SDATN ;
output EMIOPJTAGTDO ;
output EMIOPJTAGTDTN ;
output EMIOSDIO0BUSPOW ;
output EMIOSDIO0CLK ;
output EMIOSDIO0CMDO ;
output EMIOSDIO0CMDTN ;
output EMIOSDIO0LED ;
output EMIOSDIO1BUSPOW ;
output EMIOSDIO1CLK ;
output EMIOSDIO1CMDO ;
output EMIOSDIO1CMDTN ;
output EMIOSDIO1LED ;
output EMIOSPI0MO ;
output EMIOSPI0MOTN ;
output EMIOSPI0SCLKO ;
output EMIOSPI0SCLKTN ;
output EMIOSPI0SO ;
output EMIOSPI0SSNTN ;
output EMIOSPI0STN ;
output EMIOSPI1MO ;
output EMIOSPI1MOTN ;
output EMIOSPI1SCLKO ;
output EMIOSPI1SCLKTN ;
output EMIOSPI1SO ;
output EMIOSPI1SSNTN ;
output EMIOSPI1STN ;
output EMIOTRACECTL ;
output EMIOUART0DTRN ;
output EMIOUART0RTSN ;
output EMIOUART0TX ;
output EMIOUART1DTRN ;
output EMIOUART1RTSN ;
output EMIOUART1TX ;
output EMIOUSB0VBUSPWRSELECT ;
output EMIOUSB1VBUSPWRSELECT ;
output EMIOWDTRSTO ;
output EVENTEVENTO ;
output MAXIGP0ARESETN ;
output MAXIGP0ARVALID ;
output MAXIGP0AWVALID ;
output MAXIGP0BREADY ;
output MAXIGP0RREADY ;
output MAXIGP0WLAST ;
output MAXIGP0WVALID ;
output MAXIGP1ARESETN ;
output MAXIGP1ARVALID ;
output MAXIGP1AWVALID ;
output MAXIGP1BREADY ;
output MAXIGP1RREADY ;
output MAXIGP1WLAST ;
output MAXIGP1WVALID ;
output SAXIACPARESETN ;
output SAXIACPARREADY ;
output SAXIACPAWREADY ;
output SAXIACPBVALID ;
output SAXIACPRLAST ;
output SAXIACPRVALID ;
output SAXIACPWREADY ;
output SAXIGP0ARESETN ;
output SAXIGP0ARREADY ;
output SAXIGP0AWREADY ;
output SAXIGP0BVALID ;
output SAXIGP0RLAST ;
output SAXIGP0RVALID ;
output SAXIGP0WREADY ;
output SAXIGP1ARESETN ;
output SAXIGP1ARREADY ;
output SAXIGP1AWREADY ;
output SAXIGP1BVALID ;
output SAXIGP1RLAST ;
output SAXIGP1RVALID ;
output SAXIGP1WREADY ;
output SAXIHP0ARESETN ;
output SAXIHP0ARREADY ;
output SAXIHP0AWREADY ;
output SAXIHP0BVALID ;
output SAXIHP0RLAST ;
output SAXIHP0RVALID ;
output SAXIHP0WREADY ;
output SAXIHP1ARESETN ;
output SAXIHP1ARREADY ;
output SAXIHP1AWREADY ;
output SAXIHP1BVALID ;
output SAXIHP1RLAST ;
output SAXIHP1RVALID ;
output SAXIHP1WREADY ;
output SAXIHP2ARESETN ;
output SAXIHP2ARREADY ;
output SAXIHP2AWREADY ;
output SAXIHP2BVALID ;
output SAXIHP2RLAST ;
output SAXIHP2RVALID ;
output SAXIHP2WREADY ;
output SAXIHP3ARESETN ;
output SAXIHP3ARREADY ;
output SAXIHP3AWREADY ;
output SAXIHP3BVALID ;
output SAXIHP3RLAST ;
output SAXIHP3RVALID ;
output SAXIHP3WREADY ;
output [11:0] MAXIGP0ARID ;
output [11:0] MAXIGP0AWID ;
output [11:0] MAXIGP0WID ;
output [11:0] MAXIGP1ARID ;
output [11:0] MAXIGP1AWID ;
output [11:0] MAXIGP1WID ;
output [1:0] DMA0DATYPE ;
output [1:0] DMA1DATYPE ;
output [1:0] DMA2DATYPE ;
output [1:0] DMA3DATYPE ;
output [1:0] EMIOUSB0PORTINDCTL ;
output [1:0] EMIOUSB1PORTINDCTL ;
output [1:0] EVENTSTANDBYWFE ;
output [1:0] EVENTSTANDBYWFI ;
output [1:0] MAXIGP0ARBURST ;
output [1:0] MAXIGP0ARLOCK ;
output [1:0] MAXIGP0ARSIZE ;
output [1:0] MAXIGP0AWBURST ;
output [1:0] MAXIGP0AWLOCK ;
output [1:0] MAXIGP0AWSIZE ;
output [1:0] MAXIGP1ARBURST ;
output [1:0] MAXIGP1ARLOCK ;
output [1:0] MAXIGP1ARSIZE ;
output [1:0] MAXIGP1AWBURST ;
output [1:0] MAXIGP1AWLOCK ;
output [1:0] MAXIGP1AWSIZE ;
output [1:0] SAXIACPBRESP ;
output [1:0] SAXIACPRRESP ;
output [1:0] SAXIGP0BRESP ;
output [1:0] SAXIGP0RRESP ;
output [1:0] SAXIGP1BRESP ;
output [1:0] SAXIGP1RRESP ;
output [1:0] SAXIHP0BRESP ;
output [1:0] SAXIHP0RRESP ;
output [1:0] SAXIHP1BRESP ;
output [1:0] SAXIHP1RRESP ;
output [1:0] SAXIHP2BRESP ;
output [1:0] SAXIHP2RRESP ;
output [1:0] SAXIHP3BRESP ;
output [1:0] SAXIHP3RRESP ;
output [28:0] IRQP2F ;
output [2:0] EMIOSDIO0BUSVOLT ;
output [2:0] EMIOSDIO1BUSVOLT ;
output [2:0] EMIOSPI0SSON ;
output [2:0] EMIOSPI1SSON ;
output [2:0] EMIOTTC0WAVEO ;
output [2:0] EMIOTTC1WAVEO ;
output [2:0] MAXIGP0ARPROT ;
output [2:0] MAXIGP0AWPROT ;
output [2:0] MAXIGP1ARPROT ;
output [2:0] MAXIGP1AWPROT ;
output [2:0] SAXIACPBID ;
output [2:0] SAXIACPRID ;
output [2:0] SAXIHP0RACOUNT ;
output [2:0] SAXIHP1RACOUNT ;
output [2:0] SAXIHP2RACOUNT ;
output [2:0] SAXIHP3RACOUNT ;
output [31:0] EMIOTRACEDATA ;
output [31:0] FTMTP2FDEBUG ;
output [31:0] MAXIGP0ARADDR ;
output [31:0] MAXIGP0AWADDR ;
output [31:0] MAXIGP0WDATA ;
output [31:0] MAXIGP1ARADDR ;
output [31:0] MAXIGP1AWADDR ;
output [31:0] MAXIGP1WDATA ;
output [31:0] SAXIGP0RDATA ;
output [31:0] SAXIGP1RDATA ;
output [3:0] EMIOSDIO0DATAO ;
output [3:0] EMIOSDIO0DATATN ;
output [3:0] EMIOSDIO1DATAO ;
output [3:0] EMIOSDIO1DATATN ;
output [3:0] FCLKCLK ;
output [3:0] FCLKRESETN ;
output [3:0] FTMTF2PTRIGACK ;
output [3:0] FTMTP2FTRIG ;
output [3:0] MAXIGP0ARCACHE ;
output [3:0] MAXIGP0ARLEN ;
output [3:0] MAXIGP0ARQOS ;
output [3:0] MAXIGP0AWCACHE ;
output [3:0] MAXIGP0AWLEN ;
output [3:0] MAXIGP0AWQOS ;
output [3:0] MAXIGP0WSTRB ;
output [3:0] MAXIGP1ARCACHE ;
output [3:0] MAXIGP1ARLEN ;
output [3:0] MAXIGP1ARQOS ;
output [3:0] MAXIGP1AWCACHE ;
output [3:0] MAXIGP1AWLEN ;
output [3:0] MAXIGP1AWQOS ;
output [3:0] MAXIGP1WSTRB ;
output [5:0] SAXIGP0BID ;
output [5:0] SAXIGP0RID ;
output [5:0] SAXIGP1BID ;
output [5:0] SAXIGP1RID ;
output [5:0] SAXIHP0BID ;
output [5:0] SAXIHP0RID ;
output [5:0] SAXIHP0WACOUNT ;
output [5:0] SAXIHP1BID ;
output [5:0] SAXIHP1RID ;
output [5:0] SAXIHP1WACOUNT ;
output [5:0] SAXIHP2BID ;
output [5:0] SAXIHP2RID ;
output [5:0] SAXIHP2WACOUNT ;
output [5:0] SAXIHP3BID ;
output [5:0] SAXIHP3RID ;
output [5:0] SAXIHP3WACOUNT ;
output [63:0] EMIOGPIOO ;
output [63:0] EMIOGPIOTN ;
output [63:0] SAXIACPRDATA ;
output [63:0] SAXIHP0RDATA ;
output [63:0] SAXIHP1RDATA ;
output [63:0] SAXIHP2RDATA ;
output [63:0] SAXIHP3RDATA ;
output [7:0] EMIOENET0GMIITXD ;
output [7:0] EMIOENET1GMIITXD ;
output [7:0] SAXIHP0RCOUNT ;
output [7:0] SAXIHP0WCOUNT ;
output [7:0] SAXIHP1RCOUNT ;
output [7:0] SAXIHP1WCOUNT ;
output [7:0] SAXIHP2RCOUNT ;
output [7:0] SAXIHP2WCOUNT ;
output [7:0] SAXIHP3RCOUNT ;
output [7:0] SAXIHP3WCOUNT ;
inout DDRCASB ;
inout DDRCKE ;
inout DDRCKN ;
inout DDRCKP ;
inout DDRCSB ;
inout DDRDRSTB ;
inout DDRODT ;
inout DDRRASB ;
inout DDRVRN ;
inout DDRVRP ;
inout DDRWEB ;
inout PSCLK ;
inout PSPORB ;
inout PSSRSTB ;
inout [14:0] DDRA ;
inout [2:0] DDRBA ;
inout [31:0] DDRDQ ;
inout [3:0] DDRDM ;
inout [3:0] DDRDQSN ;
inout [3:0] DDRDQSP ;
inout [53:0] MIO ;
endmodule
//#### END MODULE DEFINITION FOR: PS7 ####

//#### BEGIN MODULE DEFINITION FOR :PULLDOWN ###
module PULLDOWN (O) /* synthesis syn_black_box  syn_lib_cell=1
 .noprune=1
 */;
output O /*synthesis syn_not_a_driver=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: PULLDOWN ####

//#### BEGIN MODULE DEFINITION FOR :PULLUP ###
module PULLUP (O) /* synthesis syn_black_box  syn_lib_cell=1
 .noprune=1
 */;
output O /*synthesis syn_not_a_driver=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: PULLUP ####

//#### BEGIN MODULE DEFINITION FOR :RAM128X1D ###
module RAM128X1D (DPO, SPO, A, D, DPRA, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [6:0] A ;
input [6:0] DPRA ;
input D ;
input WCLK ;
input WE ;
output DPO ;
output SPO ;
parameter INIT = 128'h0;
endmodule
//#### END MODULE DEFINITION FOR: RAM128X1D ####

//#### BEGIN MODULE DEFINITION FOR :RAM128X1S ###
module RAM128X1S (O, A0, A1, A2, A3, A4, A5, A6, D, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input A5 ;
input A6 ;
input D ;
input WCLK ;
input WE ;
output O ;
parameter INIT = 128'h00000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAM128X1S ####

//#### BEGIN MODULE DEFINITION FOR :RAM128X1S_1 ###
module RAM128X1S_1 (O, A0, A1, A2, A3, A4, A5, A6, D, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input A5 ;
input A6 ;
input D ;
input WCLK ;
input WE ;
output O ;
parameter INIT = 128'h00000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAM128X1S_1 ####

//#### BEGIN MODULE DEFINITION FOR :RAM16X1D ###
module RAM16X1D (DPO, SPO, A0, A1, A2, A3, D, DPRA0, DPRA1, DPRA2, DPRA3, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input D ;
input DPRA0 ;
input DPRA1 ;
input DPRA2 ;
input DPRA3 ;
input WCLK ;
input WE ;
output DPO ;
output SPO ;
parameter INIT = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: RAM16X1D ####

//#### BEGIN MODULE DEFINITION FOR :RAM16X1D_1 ###
module RAM16X1D_1 (DPO, SPO, A0, A1, A2, A3, D, DPRA0, DPRA1, DPRA2, DPRA3, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input D ;
input DPRA0 ;
input DPRA1 ;
input DPRA2 ;
input DPRA3 ;
input WCLK ;
input WE ;
output DPO ;
output SPO ;
parameter INIT = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: RAM16X1D_1 ####

//#### BEGIN MODULE DEFINITION FOR :RAM16X1S ###
module RAM16X1S (O, A0, A1, A2, A3, D, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input D ;
input WCLK ;
input WE ;
output O ;
parameter INIT = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: RAM16X1S ####

//#### BEGIN MODULE DEFINITION FOR :RAM16X1S_1 ###
module RAM16X1S_1 (O, A0, A1, A2, A3, D, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input D ;
input WCLK ;
input WE ;
output O ;
parameter INIT = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: RAM16X1S_1 ####

//#### BEGIN MODULE DEFINITION FOR :RAM16X2S ###
module RAM16X2S (O0, O1, A0, A1, A2, A3, D0, D1, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input D0 ;
input D1 ;
input WCLK ;
input WE ;
output O0 ;
output O1 ;
parameter INIT_00 = 16'h0000;
parameter INIT_01 = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: RAM16X2S ####

//#### BEGIN MODULE DEFINITION FOR :RAM16X4S ###
module RAM16X4S (O0, O1, O2, O3, A0, A1, A2, A3, D0, D1, D2, D3, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input D0 ;
input D1 ;
input D2 ;
input D3 ;
input WCLK ;
input WE ;
output O0 ;
output O1 ;
output O2 ;
output O3 ;
parameter INIT_00 = 16'h0000;
parameter INIT_01 = 16'h0000;
parameter INIT_02 = 16'h0000;
parameter INIT_03 = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: RAM16X4S ####

//#### BEGIN MODULE DEFINITION FOR :RAM16X8S ###
module RAM16X8S (O, A0, A1, A2, A3, D, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input WCLK ;
input WE ;
input [7:0] D ;
output [7:0] O ;
parameter INIT_00 = 16'h0000;
parameter INIT_01 = 16'h0000;
parameter INIT_02 = 16'h0000;
parameter INIT_03 = 16'h0000;
parameter INIT_04 = 16'h0000;
parameter INIT_05 = 16'h0000;
parameter INIT_06 = 16'h0000;
parameter INIT_07 = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: RAM16X8S ####

//#### BEGIN MODULE DEFINITION FOR :RAM256X1S ###
module RAM256X1S (O, A, D, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [7:0] A ;
input D ;
input WCLK ;
input WE ;
output O ;
parameter INIT = 256'h0;
endmodule
//#### END MODULE DEFINITION FOR: RAM256X1S ####

//#### BEGIN MODULE DEFINITION FOR :RAM32M ###
module RAM32M (DOA, DOB, DOC, DOD, ADDRA, ADDRB, ADDRC, ADDRD, DIA, DIB, DIC, DID, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [4:0] ADDRA ;
input [4:0] ADDRB ;
input [4:0] ADDRC ;
input [4:0] ADDRD ;
input [1:0] DIA ;
input [1:0] DIB ;
input [1:0] DIC ;
input [1:0] DID ;
input WCLK ;
input WE ;
output [1:0] DOA ;
output [1:0] DOB ;
output [1:0] DOC ;
output [1:0] DOD ;
parameter  INIT_A = 64'h0000000000000000;
parameter  INIT_B = 64'h0000000000000000;
parameter  INIT_C = 64'h0000000000000000;
parameter  INIT_D = 64'h0000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAM32M ####

//#### BEGIN MODULE DEFINITION FOR :RAM32X1D ###
module RAM32X1D (DPO, SPO, A0, A1, A2, A3, A4, D, DPRA0, DPRA1, DPRA2, DPRA3, DPRA4, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input D ;
input DPRA0 ;
input DPRA1 ;
input DPRA2 ;
input DPRA3 ;
input DPRA4 ;
input WCLK ;
input WE ;
output DPO ;
output SPO ;
parameter INIT = 32'h00000000;
endmodule
//#### END MODULE DEFINITION FOR: RAM32X1D ####

//#### BEGIN MODULE DEFINITION FOR :RAM32X1D_1 ###
module RAM32X1D_1 (DPO, SPO, A0, A1, A2, A3, A4, D, DPRA0, DPRA1, DPRA2, DPRA3, DPRA4, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input D ;
input DPRA0 ;
input DPRA1 ;
input DPRA2 ;
input DPRA3 ;
input DPRA4 ;
input WCLK ;
input WE ;
output DPO ;
output SPO ;
parameter INIT = 32'h00000000;
endmodule
//#### END MODULE DEFINITION FOR: RAM32X1D_1 ####

//#### BEGIN MODULE DEFINITION FOR :RAM32X1S ###
module RAM32X1S (O, A0, A1, A2, A3, A4, D, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input D ;
input WCLK ;
input WE ;
output O ;
parameter INIT = 32'h00000000;
endmodule
//#### END MODULE DEFINITION FOR: RAM32X1S ####

//#### BEGIN MODULE DEFINITION FOR :RAM32X1S_1 ###
module RAM32X1S_1 (O, A0, A1, A2, A3, A4, D, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input D ;
input WCLK ;
input WE ;
output O ;
parameter INIT = 32'h00000000;
endmodule
//#### END MODULE DEFINITION FOR: RAM32X1S_1 ####

//#### BEGIN MODULE DEFINITION FOR :RAM32X2S ###
module RAM32X2S (O0, O1, A0, A1, A2, A3, A4, D0, D1, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input D0 ;
input D1 ;
input WCLK ;
input WE ;
output O0 ;
output O1 ;
parameter INIT_00 = 32'h00000000;
parameter INIT_01 = 32'h00000000;
endmodule
//#### END MODULE DEFINITION FOR: RAM32X2S ####

//#### BEGIN MODULE DEFINITION FOR :RAM32X4S ###
module RAM32X4S (O0, O1, O2, O3, A0, A1, A2, A3, A4, D0, D1, D2, D3, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input D0 ;
input D1 ;
input D2 ;
input D3 ;
input WCLK ;
input WE ;
output O0 ;
output O1 ;
output O2 ;
output O3 ;
parameter INIT_00 = 32'h00000000;
parameter INIT_01 = 32'h00000000;
parameter INIT_02 = 32'h00000000;
parameter INIT_03 = 32'h00000000;
endmodule
//#### END MODULE DEFINITION FOR: RAM32X4S ####

//#### BEGIN MODULE DEFINITION FOR :RAM32X8S ###
module RAM32X8S (O, A0, A1, A2, A3, A4, D, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input WCLK ;
input WE ;
input [7:0] D ;
output [7:0] O ;
parameter INIT_00 = 32'h00000000;
parameter INIT_01 = 32'h00000000;
parameter INIT_02 = 32'h00000000;
parameter INIT_03 = 32'h00000000;
parameter INIT_04 = 32'h00000000;
parameter INIT_05 = 32'h00000000;
parameter INIT_06 = 32'h00000000;
parameter INIT_07 = 32'h00000000;
endmodule
//#### END MODULE DEFINITION FOR: RAM32X8S ####

//#### BEGIN MODULE DEFINITION FOR :RAM64M ###
module RAM64M (DOA, DOB, DOC, DOD, ADDRA, ADDRB, ADDRC, ADDRD, DIA, DIB, DIC, DID, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [5:0] ADDRA ;
input [5:0] ADDRB ;
input [5:0] ADDRC ;
input [5:0] ADDRD ;
input DIA ;
input DIB ;
input DIC ;
input DID ;
input WCLK ;
input WE ;
output DOA ;
output DOB ;
output DOC ;
output DOD ;
parameter  INIT_A = 64'h0000000000000000;
parameter  INIT_B = 64'h0000000000000000;
parameter  INIT_C = 64'h0000000000000000;
parameter  INIT_D = 64'h0000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAM64M ####

//#### BEGIN MODULE DEFINITION FOR :RAM64X1D ###
module RAM64X1D (DPO, SPO, A0, A1, A2, A3, A4, A5, D, DPRA0, DPRA1, DPRA2, DPRA3, DPRA4, DPRA5, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input A5 ;
input D ;
input DPRA0 ;
input DPRA1 ;
input DPRA2 ;
input DPRA3 ;
input DPRA4 ;
input DPRA5 ;
input WCLK ;
input WE ;
output DPO ;
output SPO ;
parameter INIT = 64'h0000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAM64X1D ####

//#### BEGIN MODULE DEFINITION FOR :RAM64X1D_1 ###
module RAM64X1D_1 (DPO, SPO, A0, A1, A2, A3, A4, A5, D, DPRA0, DPRA1, DPRA2, DPRA3, DPRA4, DPRA5, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input A5 ;
input D ;
input DPRA0 ;
input DPRA1 ;
input DPRA2 ;
input DPRA3 ;
input DPRA4 ;
input DPRA5 ;
input WCLK ;
input WE ;
output DPO ;
output SPO ;
parameter INIT = 64'h0000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAM64X1D_1 ####

//#### BEGIN MODULE DEFINITION FOR :RAM64X1S ###
module RAM64X1S (O, A0, A1, A2, A3, A4, A5, D, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input A5 ;
input D ;
input WCLK ;
input WE ;
output O ;
parameter INIT = 64'h0000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAM64X1S ####

//#### BEGIN MODULE DEFINITION FOR :RAM64X1S_1 ###
module RAM64X1S_1 (O, A0, A1, A2, A3, A4, A5, D, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input A5 ;
input D ;
input WCLK ;
input WE ;
output O ;
parameter INIT = 64'h0000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAM64X1S_1 ####

//#### BEGIN MODULE DEFINITION FOR :RAM64X2S ###
module RAM64X2S (O0, O1, A0, A1, A2, A3, A4, A5, D0, D1, WCLK, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input A5 ;
input D0 ;
input D1 ;
input WCLK ;
input WE ;
output O0 ;
output O1 ;
parameter INIT_00 = 64'h0000000000000000;
parameter INIT_01 = 64'h0000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAM64X2S ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16 ###
module RAMB16 (CASCADEOUTA, CASCADEOUTB, DOA, DOB, DOPA, DOPB, 
		 ADDRA, ADDRB, CASCADEINA, CASCADEINB, CLKA, CLKB, DIA, DIB, DIPA, DIPB, ENA, ENB, REGCEA, REGCEB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input ENA ;
input CLKA ;
input SSRA ;
input CASCADEINA ;
input REGCEA ;
input ENB ;
input CLKB ;
input SSRB ;
input CASCADEINB ;
input REGCEB ;
input [14:0] ADDRA ;
input [14:0] ADDRB ;
input [31:0] DIA ;
input [31:0] DIB ;
input [3:0] DIPA ;
input [3:0] DIPB ;
input [3:0] WEA ;
input [3:0] WEB ;
output CASCADEOUTA ;
output CASCADEOUTB ;
output [31:0] DOA ;
output [31:0] DOB ;
output [3:0] DOPA ;
output [3:0] DOPB ;
parameter DOA_REG = 0;
parameter DOB_REG = 0;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 36'h0;
parameter INIT_B = 36'h0;
parameter INIT_FILE = "NONE";
parameter INVERT_CLK_DOA_REG = "FALSE";
parameter INVERT_CLK_DOB_REG = "FALSE";
parameter RAM_EXTENSION_A = "NONE";
parameter RAM_EXTENSION_B = "NONE";
parameter READ_WIDTH_A = 0;
parameter READ_WIDTH_B = 0;
parameter SIM_COLLISION_CHECK = "ALL";
parameter SRVAL_A = 36'h0;
parameter SRVAL_B = 36'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter WRITE_WIDTH_A = 0;
parameter WRITE_WIDTH_B = 0;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16BWE ###
module RAMB16BWE (DOA, DOB, DOPA, DOPB, 
		  ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPA, DIPB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [13:0] ADDRA ;
input [13:0] ADDRB ;
input CLKA ;
input CLKB ;
input [31:0] DIA ;
input [31:0] DIB ;
input [3:0] DIPA ;
input [3:0] DIPB ;
input ENA ;
input ENB ;
input SSRA ;
input SSRB ;
input [3:0] WEA ;
input [3:0] WEB ;
output [31:0] DOA ;
output [31:0] DOB ;
output [3:0] DOPA ;
output [3:0] DOPB ;
parameter DATA_WIDTH_A = 0;
parameter DATA_WIDTH_B = 0;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 36'h0;
parameter INIT_B = 36'h0;
parameter INIT_FILE = "NONE";
parameter SIM_COLLISION_CHECK = "ALL";
parameter SRVAL_A = 36'h0;
parameter SRVAL_B = 36'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
endmodule
//#### END MODULE DEFINITION FOR: RAMB16BWE ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16BWER ###
module RAMB16BWER (DOA, DOB, DOPA, DOPB, 
		   ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPA, DIPB, ENA, ENB, REGCEA, REGCEB, RSTA, RSTB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [13:0] ADDRA ;
input [13:0] ADDRB ;
input CLKA ;
input CLKB ;
input [31:0] DIA ;
input [31:0] DIB ;
input [3:0] DIPA ;
input [3:0] DIPB ;
input ENA ;
input ENB ;
input REGCEA ;
input REGCEB ;
input RSTA ;
input RSTB ;
input [3:0] WEA ;
input [3:0] WEB ;
output [31:0] DOA ;
output [31:0] DOB ;
output [3:0] DOPA ;
output [3:0] DOPB ;
parameter DATA_WIDTH_A = 0;
parameter DATA_WIDTH_B = 0;
parameter DOA_REG = 0;
parameter DOB_REG = 0;
parameter EN_RSTRAM_A = "TRUE";
parameter EN_RSTRAM_B = "TRUE";
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 36'h0;
parameter INIT_B = 36'h0;
parameter INIT_FILE = "NONE";
parameter RSTTYPE = "SYNC";
parameter RST_PRIORITY_A = "CE";
parameter RST_PRIORITY_B = "CE";
parameter SETUP_ALL = 1000;
parameter SETUP_READ_FIRST = 3000;
parameter SIM_DEVICE = "SPARTAN3ADSP";
parameter SIM_COLLISION_CHECK = "ALL";
parameter SRVAL_A = 36'h0;
parameter SRVAL_B = 36'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
endmodule
//#### END MODULE DEFINITION FOR: RAMB16BWER ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16BWE_S18 ###
module RAMB16BWE_S18 (
	DO,
	DOP,
	ADDR,
	CLK,
	DI,
	DIP,
	EN,
	SSR,
	WE

) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLK ;
input EN ;
input SSR ;
input [1:0] WE ;
input [15:0] DI ;
input [1:0] DIP ;
input [9:0] ADDR ;
output [15:0] DO ;
output [1:0] DOP ;
parameter INIT = 18'h0;
parameter INITP_00 = 256'h0;
parameter INITP_01 = 256'h0;
parameter INITP_02 = 256'h0;
parameter INITP_03 = 256'h0;
parameter INITP_04 = 256'h0;
parameter INITP_05 = 256'h0;
parameter INITP_06 = 256'h0;
parameter INITP_07 = 256'h0;
parameter INIT_00 = 256'h0;
parameter INIT_01 = 256'h0;
parameter INIT_02 = 256'h0;
parameter INIT_03 = 256'h0;
parameter INIT_04 = 256'h0;
parameter INIT_05 = 256'h0;
parameter INIT_06 = 256'h0;
parameter INIT_07 = 256'h0;
parameter INIT_08 = 256'h0;
parameter INIT_09 = 256'h0;
parameter INIT_0A = 256'h0;
parameter INIT_0B = 256'h0;
parameter INIT_0C = 256'h0;
parameter INIT_0D = 256'h0;
parameter INIT_0E = 256'h0;
parameter INIT_0F = 256'h0;
parameter INIT_10 = 256'h0;
parameter INIT_11 = 256'h0;
parameter INIT_12 = 256'h0;
parameter INIT_13 = 256'h0;
parameter INIT_14 = 256'h0;
parameter INIT_15 = 256'h0;
parameter INIT_16 = 256'h0;
parameter INIT_17 = 256'h0;
parameter INIT_18 = 256'h0;
parameter INIT_19 = 256'h0;
parameter INIT_1A = 256'h0;
parameter INIT_1B = 256'h0;
parameter INIT_1C = 256'h0;
parameter INIT_1D = 256'h0;
parameter INIT_1E = 256'h0;
parameter INIT_1F = 256'h0;
parameter INIT_20 = 256'h0;
parameter INIT_21 = 256'h0;
parameter INIT_22 = 256'h0;
parameter INIT_23 = 256'h0;
parameter INIT_24 = 256'h0;
parameter INIT_25 = 256'h0;
parameter INIT_26 = 256'h0;
parameter INIT_27 = 256'h0;
parameter INIT_28 = 256'h0;
parameter INIT_29 = 256'h0;
parameter INIT_2A = 256'h0;
parameter INIT_2B = 256'h0;
parameter INIT_2C = 256'h0;
parameter INIT_2D = 256'h0;
parameter INIT_2E = 256'h0;
parameter INIT_2F = 256'h0;
parameter INIT_30 = 256'h0;
parameter INIT_31 = 256'h0;
parameter INIT_32 = 256'h0;
parameter INIT_33 = 256'h0;
parameter INIT_34 = 256'h0;
parameter INIT_35 = 256'h0;
parameter INIT_36 = 256'h0;
parameter INIT_37 = 256'h0;
parameter INIT_38 = 256'h0;
parameter INIT_39 = 256'h0;
parameter INIT_3A = 256'h0;
parameter INIT_3B = 256'h0;
parameter INIT_3C = 256'h0;
parameter INIT_3D = 256'h0;
parameter INIT_3E = 256'h0;
parameter INIT_3F = 256'h0;
parameter SRVAL = 18'h0;
parameter WRITE_MODE = "WRITE_FIRST";
endmodule
//#### END MODULE DEFINITION FOR: RAMB16BWE_S18 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16BWE_S18_S18 ###
module RAMB16BWE_S18_S18 (
	DOA,
	DOB,
	DOPA,
	DOPB,
	ADDRA,
	ADDRB,
	CLKA,
	CLKB,
	DIA,
	DIB,
	DIPA,
	DIPB,
	ENA,
	ENB,
	SSRA,
	SSRB,
	WEA,
	WEB

) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKA ;
input CLKB ;
input ENA ;
input ENB ;
input SSRA ;
input SSRB ;
input [1:0] WEB ;
input [1:0] WEA ;
input [15:0] DIA ;
input [15:0] DIB ;
input [1:0] DIPA ;
input [1:0] DIPB ;
input [9:0] ADDRA ;
input [9:0] ADDRB ;
output [15:0] DOA ;
output [15:0] DOB ;
output [1:0] DOPA ;
output [1:0] DOPB ;
parameter INITP_00 = 256'h0;
parameter INITP_01 = 256'h0;
parameter INITP_02 = 256'h0;
parameter INITP_03 = 256'h0;
parameter INITP_04 = 256'h0;
parameter INITP_05 = 256'h0;
parameter INITP_06 = 256'h0;
parameter INITP_07 = 256'h0;
parameter INIT_00 = 256'h0;
parameter INIT_01 = 256'h0;
parameter INIT_02 = 256'h0;
parameter INIT_03 = 256'h0;
parameter INIT_04 = 256'h0;
parameter INIT_05 = 256'h0;
parameter INIT_06 = 256'h0;
parameter INIT_07 = 256'h0;
parameter INIT_08 = 256'h0;
parameter INIT_09 = 256'h0;
parameter INIT_0A = 256'h0;
parameter INIT_0B = 256'h0;
parameter INIT_0C = 256'h0;
parameter INIT_0D = 256'h0;
parameter INIT_0E = 256'h0;
parameter INIT_0F = 256'h0;
parameter INIT_10 = 256'h0;
parameter INIT_11 = 256'h0;
parameter INIT_12 = 256'h0;
parameter INIT_13 = 256'h0;
parameter INIT_14 = 256'h0;
parameter INIT_15 = 256'h0;
parameter INIT_16 = 256'h0;
parameter INIT_17 = 256'h0;
parameter INIT_18 = 256'h0;
parameter INIT_19 = 256'h0;
parameter INIT_1A = 256'h0;
parameter INIT_1B = 256'h0;
parameter INIT_1C = 256'h0;
parameter INIT_1D = 256'h0;
parameter INIT_1E = 256'h0;
parameter INIT_1F = 256'h0;
parameter INIT_20 = 256'h0;
parameter INIT_21 = 256'h0;
parameter INIT_22 = 256'h0;
parameter INIT_23 = 256'h0;
parameter INIT_24 = 256'h0;
parameter INIT_25 = 256'h0;
parameter INIT_26 = 256'h0;
parameter INIT_27 = 256'h0;
parameter INIT_28 = 256'h0;
parameter INIT_29 = 256'h0;
parameter INIT_2A = 256'h0;
parameter INIT_2B = 256'h0;
parameter INIT_2C = 256'h0;
parameter INIT_2D = 256'h0;
parameter INIT_2E = 256'h0;
parameter INIT_2F = 256'h0;
parameter INIT_30 = 256'h0;
parameter INIT_31 = 256'h0;
parameter INIT_32 = 256'h0;
parameter INIT_33 = 256'h0;
parameter INIT_34 = 256'h0;
parameter INIT_35 = 256'h0;
parameter INIT_36 = 256'h0;
parameter INIT_37 = 256'h0;
parameter INIT_38 = 256'h0;
parameter INIT_39 = 256'h0;
parameter INIT_3A = 256'h0;
parameter INIT_3B = 256'h0;
parameter INIT_3C = 256'h0;
parameter INIT_3D = 256'h0;
parameter INIT_3E = 256'h0;
parameter INIT_3F = 256'h0;
parameter INIT_A = 18'h0;
parameter INIT_B = 18'h0;
parameter SIM_COLLISION_CHECK = "ALL";
parameter SRVAL_A = 18'h0;
parameter SRVAL_B = 18'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
endmodule
//#### END MODULE DEFINITION FOR: RAMB16BWE_S18_S18 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16BWE_S18_S9 ###
module RAMB16BWE_S18_S9 (
	DOA,
	DOB,
	DOPA,
	DOPB,
	ADDRA,
	ADDRB,
	CLKA,
	CLKB,
	DIA,
	DIB,
	DIPA,
	DIPB,
	ENA,
	ENB,
	SSRA,
	SSRB,
	WEA,
	WEB

) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [9:0] ADDRA ;
input [10:0] ADDRB ;
input CLKA ;
input CLKB ;
input [15:0] DIA ;
input [1:0] DIPA ;
input [7:0] DIB ;
input [0:0] DIPB ;
input ENA ;
input ENB ;
input SSRA ;
input SSRB ;
input [1:0] WEA ;
input WEB ;
output [15:0] DOA ;
output [1:0] DOPA ;
output [7:0] DOB ;
output [0:0] DOPB ;
parameter INITP_00 = 256'h0;
parameter INITP_01 = 256'h0;
parameter INITP_02 = 256'h0;
parameter INITP_03 = 256'h0;
parameter INITP_04 = 256'h0;
parameter INITP_05 = 256'h0;
parameter INITP_06 = 256'h0;
parameter INITP_07 = 256'h0;
parameter INIT_00 = 256'h0;
parameter INIT_01 = 256'h0;
parameter INIT_02 = 256'h0;
parameter INIT_03 = 256'h0;
parameter INIT_04 = 256'h0;
parameter INIT_05 = 256'h0;
parameter INIT_06 = 256'h0;
parameter INIT_07 = 256'h0;
parameter INIT_08 = 256'h0;
parameter INIT_09 = 256'h0;
parameter INIT_0A = 256'h0;
parameter INIT_0B = 256'h0;
parameter INIT_0C = 256'h0;
parameter INIT_0D = 256'h0;
parameter INIT_0E = 256'h0;
parameter INIT_0F = 256'h0;
parameter INIT_10 = 256'h0;
parameter INIT_11 = 256'h0;
parameter INIT_12 = 256'h0;
parameter INIT_13 = 256'h0;
parameter INIT_14 = 256'h0;
parameter INIT_15 = 256'h0;
parameter INIT_16 = 256'h0;
parameter INIT_17 = 256'h0;
parameter INIT_18 = 256'h0;
parameter INIT_19 = 256'h0;
parameter INIT_1A = 256'h0;
parameter INIT_1B = 256'h0;
parameter INIT_1C = 256'h0;
parameter INIT_1D = 256'h0;
parameter INIT_1E = 256'h0;
parameter INIT_1F = 256'h0;
parameter INIT_20 = 256'h0;
parameter INIT_21 = 256'h0;
parameter INIT_22 = 256'h0;
parameter INIT_23 = 256'h0;
parameter INIT_24 = 256'h0;
parameter INIT_25 = 256'h0;
parameter INIT_26 = 256'h0;
parameter INIT_27 = 256'h0;
parameter INIT_28 = 256'h0;
parameter INIT_29 = 256'h0;
parameter INIT_2A = 256'h0;
parameter INIT_2B = 256'h0;
parameter INIT_2C = 256'h0;
parameter INIT_2D = 256'h0;
parameter INIT_2E = 256'h0;
parameter INIT_2F = 256'h0;
parameter INIT_30 = 256'h0;
parameter INIT_31 = 256'h0;
parameter INIT_32 = 256'h0;
parameter INIT_33 = 256'h0;
parameter INIT_34 = 256'h0;
parameter INIT_35 = 256'h0;
parameter INIT_36 = 256'h0;
parameter INIT_37 = 256'h0;
parameter INIT_38 = 256'h0;
parameter INIT_39 = 256'h0;
parameter INIT_3A = 256'h0;
parameter INIT_3B = 256'h0;
parameter INIT_3C = 256'h0;
parameter INIT_3D = 256'h0;
parameter INIT_3E = 256'h0;
parameter INIT_3F = 256'h0;
parameter INIT_A = 18'h0;
parameter INIT_B = 9'h0;
parameter SIM_COLLISION_CHECK = "ALL";
parameter SRVAL_A = 18'h0;
parameter SRVAL_B = 9'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
endmodule
//#### END MODULE DEFINITION FOR: RAMB16BWE_S18_S9 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16BWE_S36 ###
module RAMB16BWE_S36 (
	DO,
	DOP,
	ADDR,
	CLK,
	DI,
	DIP,
	EN,
	SSR,
	WE

) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLK ;
input EN ;
input SSR ;
input [3:0] WE ;
input [31:0] DI ;
input [3:0] DIP ;
input [8:0] ADDR ;
output [31:0] DO ;
output [3:0] DOP ;
parameter INIT = 36'h0;
parameter INITP_00 = 256'h0;
parameter INITP_01 = 256'h0;
parameter INITP_02 = 256'h0;
parameter INITP_03 = 256'h0;
parameter INITP_04 = 256'h0;
parameter INITP_05 = 256'h0;
parameter INITP_06 = 256'h0;
parameter INITP_07 = 256'h0;
parameter INIT_00 = 256'h0;
parameter INIT_01 = 256'h0;
parameter INIT_02 = 256'h0;
parameter INIT_03 = 256'h0;
parameter INIT_04 = 256'h0;
parameter INIT_05 = 256'h0;
parameter INIT_06 = 256'h0;
parameter INIT_07 = 256'h0;
parameter INIT_08 = 256'h0;
parameter INIT_09 = 256'h0;
parameter INIT_0A = 256'h0;
parameter INIT_0B = 256'h0;
parameter INIT_0C = 256'h0;
parameter INIT_0D = 256'h0;
parameter INIT_0E = 256'h0;
parameter INIT_0F = 256'h0;
parameter INIT_10 = 256'h0;
parameter INIT_11 = 256'h0;
parameter INIT_12 = 256'h0;
parameter INIT_13 = 256'h0;
parameter INIT_14 = 256'h0;
parameter INIT_15 = 256'h0;
parameter INIT_16 = 256'h0;
parameter INIT_17 = 256'h0;
parameter INIT_18 = 256'h0;
parameter INIT_19 = 256'h0;
parameter INIT_1A = 256'h0;
parameter INIT_1B = 256'h0;
parameter INIT_1C = 256'h0;
parameter INIT_1D = 256'h0;
parameter INIT_1E = 256'h0;
parameter INIT_1F = 256'h0;
parameter INIT_20 = 256'h0;
parameter INIT_21 = 256'h0;
parameter INIT_22 = 256'h0;
parameter INIT_23 = 256'h0;
parameter INIT_24 = 256'h0;
parameter INIT_25 = 256'h0;
parameter INIT_26 = 256'h0;
parameter INIT_27 = 256'h0;
parameter INIT_28 = 256'h0;
parameter INIT_29 = 256'h0;
parameter INIT_2A = 256'h0;
parameter INIT_2B = 256'h0;
parameter INIT_2C = 256'h0;
parameter INIT_2D = 256'h0;
parameter INIT_2E = 256'h0;
parameter INIT_2F = 256'h0;
parameter INIT_30 = 256'h0;
parameter INIT_31 = 256'h0;
parameter INIT_32 = 256'h0;
parameter INIT_33 = 256'h0;
parameter INIT_34 = 256'h0;
parameter INIT_35 = 256'h0;
parameter INIT_36 = 256'h0;
parameter INIT_37 = 256'h0;
parameter INIT_38 = 256'h0;
parameter INIT_39 = 256'h0;
parameter INIT_3A = 256'h0;
parameter INIT_3B = 256'h0;
parameter INIT_3C = 256'h0;
parameter INIT_3D = 256'h0;
parameter INIT_3E = 256'h0;
parameter INIT_3F = 256'h0;
parameter SRVAL = 36'h0;
parameter WRITE_MODE = "WRITE_FIRST";
endmodule
//#### END MODULE DEFINITION FOR: RAMB16BWE_S36 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16BWE_S36_S18 ###
module RAMB16BWE_S36_S18 (
	DOA,
	DOB,
	DOPA,
	DOPB,
	ADDRA,
	ADDRB,
	CLKA,
	CLKB,
	DIA,
	DIB,
	DIPA,
	DIPB,
	ENA,
	ENB,
	SSRA,
	SSRB,
	WEA,
	WEB

) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKA ;
input CLKB ;
input ENA ;
input ENB ;
input SSRA ;
input SSRB ;
input [3:0] WEA ;
input [1:0] WEB ;
input [31:0] DIA ;
input [3:0] DIPA ;
input [15:0] DIB ;
input [1:0] DIPB ;
input [8:0] ADDRA ;
input [9:0] ADDRB ;
output [31:0] DOA ;
output [3:0] DOPA ;
output [15:0] DOB ;
output [1:0] DOPB ;
parameter INITP_00 = 256'h0;
parameter INITP_01 = 256'h0;
parameter INITP_02 = 256'h0;
parameter INITP_03 = 256'h0;
parameter INITP_04 = 256'h0;
parameter INITP_05 = 256'h0;
parameter INITP_06 = 256'h0;
parameter INITP_07 = 256'h0;
parameter INIT_00 = 256'h0;
parameter INIT_01 = 256'h0;
parameter INIT_02 = 256'h0;
parameter INIT_03 = 256'h0;
parameter INIT_04 = 256'h0;
parameter INIT_05 = 256'h0;
parameter INIT_06 = 256'h0;
parameter INIT_07 = 256'h0;
parameter INIT_08 = 256'h0;
parameter INIT_09 = 256'h0;
parameter INIT_0A = 256'h0;
parameter INIT_0B = 256'h0;
parameter INIT_0C = 256'h0;
parameter INIT_0D = 256'h0;
parameter INIT_0E = 256'h0;
parameter INIT_0F = 256'h0;
parameter INIT_10 = 256'h0;
parameter INIT_11 = 256'h0;
parameter INIT_12 = 256'h0;
parameter INIT_13 = 256'h0;
parameter INIT_14 = 256'h0;
parameter INIT_15 = 256'h0;
parameter INIT_16 = 256'h0;
parameter INIT_17 = 256'h0;
parameter INIT_18 = 256'h0;
parameter INIT_19 = 256'h0;
parameter INIT_1A = 256'h0;
parameter INIT_1B = 256'h0;
parameter INIT_1C = 256'h0;
parameter INIT_1D = 256'h0;
parameter INIT_1E = 256'h0;
parameter INIT_1F = 256'h0;
parameter INIT_20 = 256'h0;
parameter INIT_21 = 256'h0;
parameter INIT_22 = 256'h0;
parameter INIT_23 = 256'h0;
parameter INIT_24 = 256'h0;
parameter INIT_25 = 256'h0;
parameter INIT_26 = 256'h0;
parameter INIT_27 = 256'h0;
parameter INIT_28 = 256'h0;
parameter INIT_29 = 256'h0;
parameter INIT_2A = 256'h0;
parameter INIT_2B = 256'h0;
parameter INIT_2C = 256'h0;
parameter INIT_2D = 256'h0;
parameter INIT_2E = 256'h0;
parameter INIT_2F = 256'h0;
parameter INIT_30 = 256'h0;
parameter INIT_31 = 256'h0;
parameter INIT_32 = 256'h0;
parameter INIT_33 = 256'h0;
parameter INIT_34 = 256'h0;
parameter INIT_35 = 256'h0;
parameter INIT_36 = 256'h0;
parameter INIT_37 = 256'h0;
parameter INIT_38 = 256'h0;
parameter INIT_39 = 256'h0;
parameter INIT_3A = 256'h0;
parameter INIT_3B = 256'h0;
parameter INIT_3C = 256'h0;
parameter INIT_3D = 256'h0;
parameter INIT_3E = 256'h0;
parameter INIT_3F = 256'h0;
parameter INIT_A = 36'h0;
parameter INIT_B = 18'h0;
parameter SIM_COLLISION_CHECK = "ALL";
parameter SRVAL_A = 36'h0;
parameter SRVAL_B = 18'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
endmodule
//#### END MODULE DEFINITION FOR: RAMB16BWE_S36_S18 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16BWE_S36_S36 ###
module RAMB16BWE_S36_S36 (
	DOA,
	DOB,
	DOPA,
	DOPB,
	ADDRA,
	ADDRB,
	CLKA,
	CLKB,
	DIA,
	DIB,
	DIPA,
	DIPB,
	ENA,
	ENB,
	SSRA,
	SSRB,
	WEA,
	WEB

) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKA ;
input CLKB ;
input ENA ;
input ENB ;
input SSRA ;
input SSRB ;
input [3:0] WEA ;
input [3:0] WEB ;
input [31:0] DIA ;
input [31:0] DIB ;
input [3:0] DIPA ;
input [3:0] DIPB ;
input [8:0] ADDRA ;
input [8:0] ADDRB ;
output [31:0] DOA ;
output [31:0] DOB ;
output [3:0] DOPA ;
output [3:0] DOPB ;
parameter INITP_00 = 256'h0;
parameter INITP_01 = 256'h0;
parameter INITP_02 = 256'h0;
parameter INITP_03 = 256'h0;
parameter INITP_04 = 256'h0;
parameter INITP_05 = 256'h0;
parameter INITP_06 = 256'h0;
parameter INITP_07 = 256'h0;
parameter INIT_00 = 256'h0;
parameter INIT_01 = 256'h0;
parameter INIT_02 = 256'h0;
parameter INIT_03 = 256'h0;
parameter INIT_04 = 256'h0;
parameter INIT_05 = 256'h0;
parameter INIT_06 = 256'h0;
parameter INIT_07 = 256'h0;
parameter INIT_08 = 256'h0;
parameter INIT_09 = 256'h0;
parameter INIT_0A = 256'h0;
parameter INIT_0B = 256'h0;
parameter INIT_0C = 256'h0;
parameter INIT_0D = 256'h0;
parameter INIT_0E = 256'h0;
parameter INIT_0F = 256'h0;
parameter INIT_10 = 256'h0;
parameter INIT_11 = 256'h0;
parameter INIT_12 = 256'h0;
parameter INIT_13 = 256'h0;
parameter INIT_14 = 256'h0;
parameter INIT_15 = 256'h0;
parameter INIT_16 = 256'h0;
parameter INIT_17 = 256'h0;
parameter INIT_18 = 256'h0;
parameter INIT_19 = 256'h0;
parameter INIT_1A = 256'h0;
parameter INIT_1B = 256'h0;
parameter INIT_1C = 256'h0;
parameter INIT_1D = 256'h0;
parameter INIT_1E = 256'h0;
parameter INIT_1F = 256'h0;
parameter INIT_20 = 256'h0;
parameter INIT_21 = 256'h0;
parameter INIT_22 = 256'h0;
parameter INIT_23 = 256'h0;
parameter INIT_24 = 256'h0;
parameter INIT_25 = 256'h0;
parameter INIT_26 = 256'h0;
parameter INIT_27 = 256'h0;
parameter INIT_28 = 256'h0;
parameter INIT_29 = 256'h0;
parameter INIT_2A = 256'h0;
parameter INIT_2B = 256'h0;
parameter INIT_2C = 256'h0;
parameter INIT_2D = 256'h0;
parameter INIT_2E = 256'h0;
parameter INIT_2F = 256'h0;
parameter INIT_30 = 256'h0;
parameter INIT_31 = 256'h0;
parameter INIT_32 = 256'h0;
parameter INIT_33 = 256'h0;
parameter INIT_34 = 256'h0;
parameter INIT_35 = 256'h0;
parameter INIT_36 = 256'h0;
parameter INIT_37 = 256'h0;
parameter INIT_38 = 256'h0;
parameter INIT_39 = 256'h0;
parameter INIT_3A = 256'h0;
parameter INIT_3B = 256'h0;
parameter INIT_3C = 256'h0;
parameter INIT_3D = 256'h0;
parameter INIT_3E = 256'h0;
parameter INIT_3F = 256'h0;
parameter INIT_A = 36'h0;
parameter INIT_B = 36'h0;
parameter SIM_COLLISION_CHECK = "ALL";
parameter SRVAL_A = 36'h0;
parameter SRVAL_B = 36'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
endmodule
//#### END MODULE DEFINITION FOR: RAMB16BWE_S36_S36 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16BWE_S36_S9 ###
module RAMB16BWE_S36_S9 (
	DOA,
	DOB,
	DOPA,
	DOPB,
	ADDRA,
	ADDRB,
	CLKA,
	CLKB,
	DIA,
	DIB,
	DIPA,
	DIPB,
	ENA,
	ENB,
	SSRA,
	SSRB,
	WEA,
	WEB

) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [8:0]  ADDRA ;
input [10:0] ADDRB ;
input CLKA ;
input CLKB ;
input ENA ;
input ENB ;
input SSRA ;
input SSRB ;
input [3:0] WEA ;
input WEB ;
input [31:0] DIA ;
input [3:0] DIPA ;
input [7:0] DIB ;
input [0:0] DIPB ;
output [31:0] DOA ;
output [3:0]  DOPA ;
output [7:0]  DOB ;
output [0:0]  DOPB ;
parameter INITP_00 = 256'h0;
parameter INITP_01 = 256'h0;
parameter INITP_02 = 256'h0;
parameter INITP_03 = 256'h0;
parameter INITP_04 = 256'h0;
parameter INITP_05 = 256'h0;
parameter INITP_06 = 256'h0;
parameter INITP_07 = 256'h0;
parameter INIT_00 = 256'h0;
parameter INIT_01 = 256'h0;
parameter INIT_02 = 256'h0;
parameter INIT_03 = 256'h0;
parameter INIT_04 = 256'h0;
parameter INIT_05 = 256'h0;
parameter INIT_06 = 256'h0;
parameter INIT_07 = 256'h0;
parameter INIT_08 = 256'h0;
parameter INIT_09 = 256'h0;
parameter INIT_0A = 256'h0;
parameter INIT_0B = 256'h0;
parameter INIT_0C = 256'h0;
parameter INIT_0D = 256'h0;
parameter INIT_0E = 256'h0;
parameter INIT_0F = 256'h0;
parameter INIT_10 = 256'h0;
parameter INIT_11 = 256'h0;
parameter INIT_12 = 256'h0;
parameter INIT_13 = 256'h0;
parameter INIT_14 = 256'h0;
parameter INIT_15 = 256'h0;
parameter INIT_16 = 256'h0;
parameter INIT_17 = 256'h0;
parameter INIT_18 = 256'h0;
parameter INIT_19 = 256'h0;
parameter INIT_1A = 256'h0;
parameter INIT_1B = 256'h0;
parameter INIT_1C = 256'h0;
parameter INIT_1D = 256'h0;
parameter INIT_1E = 256'h0;
parameter INIT_1F = 256'h0;
parameter INIT_20 = 256'h0;
parameter INIT_21 = 256'h0;
parameter INIT_22 = 256'h0;
parameter INIT_23 = 256'h0;
parameter INIT_24 = 256'h0;
parameter INIT_25 = 256'h0;
parameter INIT_26 = 256'h0;
parameter INIT_27 = 256'h0;
parameter INIT_28 = 256'h0;
parameter INIT_29 = 256'h0;
parameter INIT_2A = 256'h0;
parameter INIT_2B = 256'h0;
parameter INIT_2C = 256'h0;
parameter INIT_2D = 256'h0;
parameter INIT_2E = 256'h0;
parameter INIT_2F = 256'h0;
parameter INIT_30 = 256'h0;
parameter INIT_31 = 256'h0;
parameter INIT_32 = 256'h0;
parameter INIT_33 = 256'h0;
parameter INIT_34 = 256'h0;
parameter INIT_35 = 256'h0;
parameter INIT_36 = 256'h0;
parameter INIT_37 = 256'h0;
parameter INIT_38 = 256'h0;
parameter INIT_39 = 256'h0;
parameter INIT_3A = 256'h0;
parameter INIT_3B = 256'h0;
parameter INIT_3C = 256'h0;
parameter INIT_3D = 256'h0;
parameter INIT_3E = 256'h0;
parameter INIT_3F = 256'h0;
parameter INIT_A = 36'h0;
parameter INIT_B = 9'h0;
parameter SIM_COLLISION_CHECK = "ALL";
parameter SRVAL_A = 36'h0;
parameter SRVAL_B = 9'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
endmodule
//#### END MODULE DEFINITION FOR: RAMB16BWE_S36_S9 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S1 ###
module RAMB16_S1 (DO, ADDR, CLK, DI, EN, SSR, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [13:0] ADDR ;
input [0:0] DI ;
input EN ;
input CLK ;
input WE ;
input SSR ;
output [0:0] DO ;
parameter INIT = 1'h0;
parameter SRVAL = 1'h0;
parameter WRITE_MODE = "WRITE_FIRST";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S1 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S18 ###
module RAMB16_S18 (DO, DOP, ADDR, CLK, DI, DIP, EN, SSR, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [9:0] ADDR ;
input [15:0] DI ;
input [1:0] DIP ;
input EN ;
input CLK ;
input WE ;
input SSR ;
output [15:0] DO ;
output [1:0] DOP ;
parameter INIT = 18'h0;
parameter SRVAL = 18'h0;
parameter WRITE_MODE = "WRITE_FIRST";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S18 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S18_S18 ###
module RAMB16_S18_S18 (DOA, DOB, DOPA, DOPB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPA, DIPB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [9:0] ADDRA ;
input [15:0] DIA ;
input [1:0] DIPA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [9:0] ADDRB ;
input [15:0] DIB ;
input [1:0] DIPB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [15:0] DOA ;
output [1:0] DOPA ;
output [15:0] DOB ;
output [1:0] DOPB ;
parameter INIT_A = 18'h0;
parameter INIT_B = 18'h0;
parameter SRVAL_A = 18'h0;
parameter SRVAL_B = 18'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S18_S18 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S18_S36 ###
module RAMB16_S18_S36 (DOA, DOB, DOPA, DOPB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPA, DIPB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [9:0] ADDRA ;
input [15:0] DIA ;
input [1:0] DIPA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [8:0] ADDRB ;
input [31:0] DIB ;
input [3:0] DIPB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [15:0] DOA ;
output [1:0] DOPA ;
output [31:0] DOB ;
output [3:0] DOPB ;
parameter INIT_A = 18'h0;
parameter INIT_B = 36'h0;
parameter SRVAL_A = 18'h0;
parameter SRVAL_B = 36'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S18_S36 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S1_S1 ###
module RAMB16_S1_S1 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [13:0] ADDRA ;
input [0:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [13:0] ADDRB ;
input [0:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [0:0] DOA ;
output [0:0] DOB ;
parameter INIT_A = 1'h0;
parameter INIT_B = 1'h0;
parameter SRVAL_A = 1'h0;
parameter SRVAL_B = 1'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S1_S1 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S1_S18 ###
module RAMB16_S1_S18 (DOA, DOB, DOPB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [13:0] ADDRA ;
input [0:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [9:0] ADDRB ;
input [15:0] DIB ;
input [1:0] DIPB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [0:0] DOA ;
output [15:0] DOB ;
output [1:0] DOPB ;
parameter INIT_A = 1'h0;
parameter INIT_B = 18'h0;
parameter SRVAL_A = 1'h0;
parameter SRVAL_B = 18'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S1_S18 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S1_S2 ###
module RAMB16_S1_S2 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [13:0] ADDRA ;
input [0:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [12:0] ADDRB ;
input [1:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [0:0] DOA ;
output [1:0] DOB ;
parameter INIT_A = 1'h0;
parameter INIT_B = 2'h0;
parameter SRVAL_A = 1'h0;
parameter SRVAL_B = 2'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S1_S2 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S1_S36 ###
module RAMB16_S1_S36 (DOA, DOB, DOPB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [13:0] ADDRA ;
input [0:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [8:0] ADDRB ;
input [31:0] DIB ;
input [3:0] DIPB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [0:0] DOA ;
output [31:0] DOB ;
output [3:0] DOPB ;
parameter INIT_A = 1'h0;
parameter INIT_B = 36'h0;
parameter SRVAL_A = 1'h0;
parameter SRVAL_B = 36'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S1_S36 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S1_S4 ###
module RAMB16_S1_S4 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [13:0] ADDRA ;
input [0:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [11:0] ADDRB ;
input [3:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [0:0] DOA ;
output [3:0] DOB ;
parameter INIT_A = 1'h0;
parameter INIT_B = 4'h0;
parameter SRVAL_A = 1'h0;
parameter SRVAL_B = 4'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S1_S4 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S1_S9 ###
module RAMB16_S1_S9 (DOA, DOB, DOPB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [13:0] ADDRA ;
input [0:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [10:0] ADDRB ;
input [7:0] DIB ;
input [0:0] DIPB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [0:0] DOA ;
output [7:0] DOB ;
output [0:0] DOPB ;
parameter INIT_A = 1'h0;
parameter INIT_B = 9'h0;
parameter SRVAL_A = 1'h0;
parameter SRVAL_B = 9'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S1_S9 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S2 ###
module RAMB16_S2 (DO, ADDR, CLK, DI, EN, SSR, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [12:0] ADDR ;
input [1:0] DI ;
input EN ;
input CLK ;
input WE ;
input SSR ;
output [1:0] DO ;
parameter INIT = 2'h0;
parameter SRVAL = 2'h0;
parameter WRITE_MODE = "WRITE_FIRST";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S2 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S2_S18 ###
module RAMB16_S2_S18 (DOA, DOB, DOPB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [12:0] ADDRA ;
input [1:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [9:0] ADDRB ;
input [15:0] DIB ;
input [1:0] DIPB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [1:0] DOA ;
output [15:0] DOB ;
output [1:0] DOPB ;
parameter INIT_A = 2'h0;
parameter INIT_B = 18'h0;
parameter SRVAL_A = 2'h0;
parameter SRVAL_B = 18'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S2_S18 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S2_S2 ###
module RAMB16_S2_S2 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [12:0] ADDRA ;
input [1:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [12:0] ADDRB ;
input [1:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [1:0] DOA ;
output [1:0] DOB ;
parameter INIT_A = 2'h0;
parameter INIT_B = 2'h0;
parameter SRVAL_A = 2'h0;
parameter SRVAL_B = 2'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S2_S2 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S2_S36 ###
module RAMB16_S2_S36 (DOA, DOB, DOPB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [12:0] ADDRA ;
input [1:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [8:0] ADDRB ;
input [31:0] DIB ;
input [3:0] DIPB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [1:0] DOA ;
output [31:0] DOB ;
output [3:0] DOPB ;
parameter INIT_A = 2'h0;
parameter INIT_B = 36'h0;
parameter SRVAL_A = 2'h0;
parameter SRVAL_B = 36'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S2_S36 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S2_S4 ###
module RAMB16_S2_S4 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [12:0] ADDRA ;
input [1:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [11:0] ADDRB ;
input [3:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [1:0] DOA ;
output [3:0] DOB ;
parameter INIT_A = 2'h0;
parameter INIT_B = 4'h0;
parameter SRVAL_A = 2'h0;
parameter SRVAL_B = 4'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S2_S4 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S2_S9 ###
module RAMB16_S2_S9 (DOA, DOB, DOPB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [12:0] ADDRA ;
input [1:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [10:0] ADDRB ;
input [7:0] DIB ;
input [0:0] DIPB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [1:0] DOA ;
output [7:0] DOB ;
output [0:0] DOPB ;
parameter INIT_A = 2'h0;
parameter INIT_B = 9'h0;
parameter SRVAL_A = 2'h0;
parameter SRVAL_B = 9'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S2_S9 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S36 ###
module RAMB16_S36 (DO, DOP, ADDR, CLK, DI, DIP, EN, SSR, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [8:0] ADDR ;
input [31:0] DI ;
input [3:0] DIP ;
input EN ;
input CLK ;
input WE ;
input SSR ;
output [31:0] DO ;
output [3:0] DOP ;
parameter INIT = 36'h0;
parameter SRVAL = 36'h0;
parameter WRITE_MODE = "WRITE_FIRST";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S36 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S36_S36 ###
module RAMB16_S36_S36 (DOA, DOB, DOPA, DOPB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPA, DIPB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [8:0] ADDRA ;
input [31:0] DIA ;
input [3:0] DIPA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [8:0] ADDRB ;
input [31:0] DIB ;
input [3:0] DIPB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [31:0] DOA ;
output [3:0] DOPA ;
output [31:0] DOB ;
output [3:0] DOPB ;
parameter INIT_A = 36'h0;
parameter INIT_B = 36'h0;
parameter SRVAL_A = 36'h0;
parameter SRVAL_B = 36'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S36_S36 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S4 ###
module RAMB16_S4 (DO, ADDR, CLK, DI, EN, SSR, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [11:0] ADDR ;
input [3:0] DI ;
input EN ;
input CLK ;
input WE ;
input SSR ;
output [3:0] DO ;
parameter INIT = 4'h0;
parameter SRVAL = 4'h0;
parameter WRITE_MODE = "WRITE_FIRST";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S4 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S4_S18 ###
module RAMB16_S4_S18 (DOA, DOB, DOPB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [11:0] ADDRA ;
input [3:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [9:0] ADDRB ;
input [15:0] DIB ;
input [1:0] DIPB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [3:0] DOA ;
output [15:0] DOB ;
output [1:0] DOPB ;
parameter INIT_A = 4'h0;
parameter INIT_B = 18'h0;
parameter SRVAL_A = 4'h0;
parameter SRVAL_B = 18'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S4_S18 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S4_S36 ###
module RAMB16_S4_S36 (DOA, DOB, DOPB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [11:0] ADDRA ;
input [3:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [8:0] ADDRB ;
input [31:0] DIB ;
input [3:0] DIPB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [3:0] DOA ;
output [31:0] DOB ;
output [3:0] DOPB ;
parameter INIT_A = 4'h0;
parameter INIT_B = 36'h0;
parameter SRVAL_A = 4'h0;
parameter SRVAL_B = 36'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S4_S36 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S4_S4 ###
module RAMB16_S4_S4 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [11:0] ADDRA ;
input [3:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [11:0] ADDRB ;
input [3:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [3:0] DOA ;
output [3:0] DOB ;
parameter INIT_A = 4'h0;
parameter INIT_B = 4'h0;
parameter SRVAL_A = 4'h0;
parameter SRVAL_B = 4'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S4_S4 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S4_S9 ###
module RAMB16_S4_S9 (DOA, DOB, DOPB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [11:0] ADDRA ;
input [3:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [10:0] ADDRB ;
input [7:0] DIB ;
input [0:0] DIPB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [3:0] DOA ;
output [7:0] DOB ;
output [0:0] DOPB ;
parameter INIT_A = 4'h0;
parameter INIT_B = 9'h0;
parameter SRVAL_A = 4'h0;
parameter SRVAL_B = 9'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S4_S9 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S9 ###
module RAMB16_S9 (DO, DOP, ADDR, CLK, DI, DIP, EN, SSR, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [10:0] ADDR ;
input [7:0] DI ;
input [0:0] DIP ;
input EN ;
input CLK ;
input WE ;
input SSR ;
output [7:0] DO ;
output [0:0] DOP ;
parameter INIT = 9'h0;
parameter SRVAL = 9'h0;
parameter WRITE_MODE = "WRITE_FIRST";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S9 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S9_S18 ###
module RAMB16_S9_S18 (DOA, DOB, DOPA, DOPB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPA, DIPB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [10:0] ADDRA ;
input [7:0] DIA ;
input [0:0] DIPA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [9:0] ADDRB ;
input [15:0] DIB ;
input [1:0] DIPB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [7:0] DOA ;
output [0:0] DOPA ;
output [15:0] DOB ;
output [1:0] DOPB ;
parameter INIT_A = 9'h0;
parameter INIT_B = 18'h0;
parameter SRVAL_A = 9'h0;
parameter SRVAL_B = 18'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S9_S18 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S9_S36 ###
module RAMB16_S9_S36 (DOA, DOB, DOPA, DOPB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPA, DIPB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [10:0] ADDRA ;
input [7:0] DIA ;
input [0:0] DIPA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [8:0] ADDRB ;
input [31:0] DIB ;
input [3:0] DIPB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [7:0] DOA ;
output [0:0] DOPA ;
output [31:0] DOB ;
output [3:0] DOPB ;
parameter INIT_A = 9'h0;
parameter INIT_B = 36'h0;
parameter SRVAL_A = 9'h0;
parameter SRVAL_B = 36'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S9_S36 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB16_S9_S9 ###
module RAMB16_S9_S9 (DOA, DOB, DOPA, DOPB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPA, DIPB, ENA, ENB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [10:0] ADDRA ;
input [7:0] DIA ;
input [0:0] DIPA ;
input ENA ;
input CLKA ;
input WEA ;
input SSRA ;
input [10:0] ADDRB ;
input [7:0] DIB ;
input [0:0] DIPB ;
input ENB ;
input CLKB ;
input WEB ;
input SSRB ;
output [7:0] DOA ;
output [0:0] DOPA ;
output [7:0] DOB ;
output [0:0] DOPB ;
parameter INIT_A = 9'h0;
parameter INIT_B = 9'h0;
parameter SRVAL_A = 9'h0;
parameter SRVAL_B = 9'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB16_S9_S9 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB18 ###
module RAMB18 (DOA, DOB, DOPA, DOPB,
	       ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, DIPA, DIPB, ENA, ENB, REGCEA, REGCEB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input ENA ;
input CLKA ;
input SSRA ;
input REGCEA ;
input ENB ;
input CLKB ;
input SSRB ;
input REGCEB ;
input [13:0] ADDRA ;
input [13:0] ADDRB ;
input [15:0] DIA ;
input [15:0] DIB ;
input [1:0] DIPA ;
input [1:0] DIPB ;
input [1:0] WEA ;
input [1:0] WEB ;
output [15:0] DOA ;
output [15:0] DOB ;
output [1:0] DOPA ;
output [1:0] DOPB ;
parameter DOA_REG = 0;
parameter DOB_REG = 0;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 18'h0;
parameter INIT_B = 18'h0;
parameter INIT_FILE = "NONE";
parameter READ_WIDTH_A = 0;
parameter READ_WIDTH_B = 0;
parameter SIM_COLLISION_CHECK = "ALL";
parameter SIM_MODE = "SAFE";
parameter SRVAL_A = 18'h0;
parameter SRVAL_B = 18'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter WRITE_WIDTH_A = 0;
parameter WRITE_WIDTH_B = 0;
endmodule
//#### END MODULE DEFINITION FOR: RAMB18 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB18E1 ###
module RAMB18E1 (DOADO, DOBDO, DOPADOP, DOPBDOP,
		 ADDRARDADDR, ADDRBWRADDR, CLKARDCLK, CLKBWRCLK, DIADI, DIBDI, DIPADIP, DIPBDIP, ENARDEN, ENBWREN, REGCEAREGCE, REGCEB, RSTRAMARSTRAM, RSTRAMB, RSTREGARSTREG, RSTREGB, WEA, WEBWE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLKARDCLK ;
input CLKBWRCLK ;
input ENARDEN ;
input ENBWREN ;
input REGCEAREGCE ;
input REGCEB ;
input RSTRAMARSTRAM ;
input RSTRAMB ;
input RSTREGARSTREG ;
input RSTREGB ;
input [13:0] ADDRARDADDR ;
input [13:0] ADDRBWRADDR ;
input [15:0] DIADI ;
input [15:0] DIBDI ;
input [1:0] DIPADIP ;
input [1:0] DIPBDIP ;
input [1:0] WEA ;
input [3:0] WEBWE ;
output [15:0] DOADO ;
output [15:0] DOBDO ;
output [1:0] DOPADOP ;
output [1:0] DOPBDOP ;
parameter DOA_REG = 0;
parameter DOB_REG = 0;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 18'h0;
parameter INIT_B = 18'h0;
parameter INIT_FILE = "NONE";
parameter RAM_MODE = "TDP";
parameter RDADDR_COLLISION_HWCONFIG = "DELAYED_WRITE";
parameter READ_WIDTH_A = 0;
parameter READ_WIDTH_B = 0;
parameter RSTREG_PRIORITY_A = "RSTREG";
parameter RSTREG_PRIORITY_B = "RSTREG";
parameter SIM_COLLISION_CHECK = "ALL";
parameter SIM_DEVICE = "VIRTEX6";
parameter SRVAL_A = 18'h0;
parameter SRVAL_B = 18'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter WRITE_WIDTH_A = 0;
parameter WRITE_WIDTH_B = 0;
endmodule
//#### END MODULE DEFINITION FOR: RAMB18E1 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB18SDP ###
module RAMB18SDP (DO, DOP, 
		  DI, DIP, RDADDR, RDCLK, RDEN, REGCE, SSR, WE, WRADDR, WRCLK, WREN) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input RDCLK ;
input RDEN ;
input REGCE ;
input SSR ;
input WRCLK ;
input WREN ;
input [8:0] WRADDR ;
input [8:0] RDADDR ;
input [31:0] DI ;
input [3:0] DIP ;
input [3:0] WE ;
output [31:0] DO ;
output [3:0] DOP ;
parameter DO_REG = 0;
parameter INIT = 36'h0;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_FILE = "NONE";
parameter SIM_COLLISION_CHECK = "ALL";
parameter SIM_MODE = "SAFE";
parameter SRVAL = 36'h0;
endmodule
//#### END MODULE DEFINITION FOR: RAMB18SDP ####

//#### BEGIN MODULE DEFINITION FOR :RAMB32_S64_ECC ###
module RAMB32_S64_ECC (
 DO,
 STATUS,

 DI,
 RDADDR,
 RDCLK,
 RDEN,
 SSR,
 WRADDR,
 WRCLK,
 WREN
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input RDCLK ;
input RDEN ;
input SSR ;
input WRCLK ;
input WREN ;
input [63:0] DI ;
input [8:0]  RDADDR ;
input [8:0]  WRADDR ;
output [1:0] STATUS ;
output [63:0] DO ;
parameter DO_REG = 0;
parameter SIM_COLLISION_CHECK = "ALL";
endmodule
//#### END MODULE DEFINITION FOR: RAMB32_S64_ECC ####

//#### BEGIN MODULE DEFINITION FOR :RAMB36 ###
module RAMB36 (CASCADEOUTLATA, CASCADEOUTLATB, CASCADEOUTREGA, CASCADEOUTREGB, DOA, DOB, DOPA, DOPB,
	       ADDRA, ADDRB, CASCADEINLATA, CASCADEINLATB, CASCADEINREGA, CASCADEINREGB, CLKA, CLKB, DIA, DIB, DIPA, DIPB, ENA, ENB, REGCEA, REGCEB, SSRA, SSRB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input ENA ;
input CLKA ;
input SSRA ;
input CASCADEINLATA ;
input CASCADEINREGA ;
input REGCEA ;
input ENB ;
input CLKB ;
input SSRB ;
input CASCADEINLATB ;
input CASCADEINREGB ;
input REGCEB ;
input [15:0] ADDRA ;
input [15:0] ADDRB ;
input [31:0] DIA ;
input [31:0] DIB ;
input [3:0] DIPA ;
input [3:0] DIPB ;
input [3:0] WEA ;
input [3:0] WEB ;
output CASCADEOUTLATA ;
output CASCADEOUTREGA ;
output CASCADEOUTLATB ;
output CASCADEOUTREGB ;
output [31:0] DOA ;
output [31:0] DOB ;
output [3:0] DOPA ;
output [3:0] DOPB ;
parameter DOA_REG = 0;
parameter DOB_REG = 0;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_40 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_41 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_42 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_43 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_44 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_45 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_46 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_47 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_48 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_49 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_50 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_51 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_52 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_53 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_54 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_55 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_56 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_57 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_58 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_59 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_60 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_61 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_62 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_63 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_64 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_65 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_66 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_67 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_68 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_69 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_70 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_71 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_72 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_73 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_74 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_75 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_76 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_77 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_78 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_79 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 36'h0;
parameter INIT_B = 36'h0;
parameter INIT_FILE = "NONE";
parameter RAM_EXTENSION_A = "NONE";
parameter RAM_EXTENSION_B = "NONE";
parameter READ_WIDTH_A = 0;
parameter READ_WIDTH_B = 0;
parameter SIM_COLLISION_CHECK = "ALL";
parameter SIM_MODE = "SAFE";
parameter SRVAL_A = 36'h0;
parameter SRVAL_B = 36'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter WRITE_WIDTH_A = 0;
parameter WRITE_WIDTH_B = 0;
endmodule
//#### END MODULE DEFINITION FOR: RAMB36 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB36E1 ###
module RAMB36E1 (CASCADEOUTA, CASCADEOUTB, DBITERR, DOADO, DOBDO, DOPADOP, DOPBDOP, ECCPARITY, RDADDRECC, SBITERR, 
		 ADDRARDADDR, ADDRBWRADDR, CASCADEINA, CASCADEINB, CLKARDCLK, CLKBWRCLK, DIADI, DIBDI, DIPADIP, DIPBDIP, ENARDEN, ENBWREN, INJECTDBITERR, INJECTSBITERR, REGCEAREGCE, REGCEB, RSTRAMARSTRAM, RSTRAMB, RSTREGARSTREG, RSTREGB, WEA, WEBWE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input ENARDEN ;
input CLKARDCLK ;
input RSTRAMARSTRAM ;
input RSTREGARSTREG ;
input CASCADEINA ;
input REGCEAREGCE ;
input ENBWREN ;
input CLKBWRCLK ;
input RSTRAMB ;
input RSTREGB ;
input CASCADEINB ;
input REGCEB ;
input INJECTDBITERR ;
input INJECTSBITERR ;
input [15:0] ADDRARDADDR ;
input [15:0] ADDRBWRADDR ;
input [31:0] DIADI ;
input [31:0] DIBDI ;
input [3:0] DIPADIP ;
input [3:0] DIPBDIP ;
input [3:0] WEA ;
input [7:0] WEBWE ;
output CASCADEOUTA ;
output CASCADEOUTB ;
output [31:0] DOADO ;
output [31:0] DOBDO ;
output [3:0] DOPADOP ;
output [3:0] DOPBDOP ;
output [7:0] ECCPARITY ;
output [8:0] RDADDRECC ;
output SBITERR ;
output DBITERR ;
parameter DOA_REG = 0;
parameter DOB_REG = 0;
parameter EN_ECC_READ = "FALSE";
parameter EN_ECC_WRITE = "FALSE";
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_40 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_41 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_42 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_43 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_44 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_45 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_46 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_47 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_48 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_49 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_50 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_51 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_52 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_53 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_54 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_55 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_56 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_57 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_58 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_59 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_60 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_61 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_62 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_63 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_64 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_65 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_66 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_67 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_68 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_69 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_70 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_71 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_72 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_73 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_74 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_75 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_76 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_77 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_78 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_79 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 36'h0;
parameter INIT_B = 36'h0;
parameter INIT_FILE = "NONE";
parameter RAM_EXTENSION_A = "NONE";
parameter RAM_EXTENSION_B = "NONE";
parameter RAM_MODE = "TDP";
parameter RDADDR_COLLISION_HWCONFIG = "DELAYED_WRITE";
parameter READ_WIDTH_A = 0;
parameter READ_WIDTH_B = 0;
parameter RSTREG_PRIORITY_A = "RSTREG";
parameter RSTREG_PRIORITY_B = "RSTREG";
parameter SIM_COLLISION_CHECK = "ALL";
parameter SIM_DEVICE = "VIRTEX6";
parameter SRVAL_A = 36'h0;
parameter SRVAL_B = 36'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter WRITE_WIDTH_A = 0;
parameter WRITE_WIDTH_B = 0;
endmodule
//#### END MODULE DEFINITION FOR: RAMB36E1 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB36SDP ###
module RAMB36SDP (DBITERR, DO, DOP, ECCPARITY, SBITERR, 
		  DI, DIP, RDADDR, RDCLK, RDEN, REGCE, SSR, WE, WRADDR, WRCLK, WREN) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input RDCLK ;
input RDEN ;
input REGCE ;
input SSR ;
input WRCLK ;
input WREN ;
input [8:0] WRADDR ;
input [8:0] RDADDR ;
input [63:0] DI ;
input [7:0] DIP ;
input [7:0] WE ;
output DBITERR ;
output SBITERR ;
output [63:0] DO ;
output [7:0] DOP ;
output [7:0] ECCPARITY ;
parameter DO_REG = 0;
parameter EN_ECC_READ = "FALSE";
parameter EN_ECC_SCRUB = "FALSE";
parameter EN_ECC_WRITE = "FALSE";
parameter INIT = 72'h0;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_40 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_41 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_42 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_43 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_44 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_45 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_46 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_47 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_48 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_49 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_50 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_51 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_52 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_53 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_54 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_55 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_56 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_57 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_58 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_59 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_60 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_61 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_62 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_63 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_64 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_65 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_66 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_67 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_68 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_69 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_70 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_71 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_72 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_73 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_74 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_75 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_76 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_77 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_78 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_79 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_FILE = "NONE";
parameter SIM_COLLISION_CHECK = "ALL";
parameter SIM_MODE = "SAFE";
parameter SRVAL = 72'h0;
endmodule
//#### END MODULE DEFINITION FOR: RAMB36SDP ####

//#### BEGIN MODULE DEFINITION FOR :RAMB36SDP_EXP ###
module RAMB36SDP_EXP (DBITERR, DO, DOP, ECCPARITY, SBITERR, 
		      DI, DIP, RDADDRL, RDADDRU, RDCLKL, RDCLKU, RDENL, RDENU, RDRCLKL, RDRCLKU, REGCEL, REGCEU, SSRL, SSRU, WEL, WEU, WRADDRL, WRADDRU, WRCLKL, WRCLKU, WRENL, WRENU ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input RDCLKL ;
input RDCLKU ;
input RDENL ;
input RDENU ;
input RDRCLKL ;
input RDRCLKU ;
input REGCEL ;
input REGCEU ;
input SSRL ;
input SSRU ;
input WRCLKL ;
input WRCLKU ;
input WRENL ;
input WRENU ;
input [14:0] RDADDRU ;
input [14:0] WRADDRU ;
input [15:0] RDADDRL ;
input [15:0] WRADDRL ;
input [63:0] DI ;
input [7:0] DIP ;
input [7:0] WEL ;
input [7:0] WEU ;
output DBITERR ;
output SBITERR ;
output [63:0] DO ;
output [7:0] DOP ;
output [7:0] ECCPARITY ;
parameter DO_REG = 0;
parameter EN_ECC_READ = "FALSE";
parameter EN_ECC_SCRUB = "FALSE";
parameter EN_ECC_WRITE = "FALSE";
parameter INIT = 72'h0;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_40 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_41 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_42 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_43 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_44 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_45 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_46 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_47 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_48 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_49 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_50 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_51 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_52 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_53 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_54 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_55 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_56 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_57 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_58 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_59 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_60 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_61 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_62 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_63 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_64 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_65 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_66 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_67 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_68 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_69 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_70 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_71 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_72 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_73 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_74 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_75 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_76 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_77 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_78 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_79 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_FILE = "NONE";
parameter SIM_COLLISION_CHECK = "ALL";
parameter SIM_MODE = "SAFE";
parameter SRVAL = 72'h0;
endmodule
//#### END MODULE DEFINITION FOR: RAMB36SDP_EXP ####

//#### BEGIN MODULE DEFINITION FOR :RAMB36_EXP ###
module RAMB36_EXP (CASCADEOUTLATA, CASCADEOUTLATB, CASCADEOUTREGA, CASCADEOUTREGB, DOA, DOB, DOPA, DOPB,
		   ADDRAL, ADDRAU, ADDRBL, ADDRBU, CASCADEINLATA, CASCADEINLATB, CASCADEINREGA, CASCADEINREGB, CLKAL, CLKAU, CLKBL, CLKBU, DIA, DIB, DIPA, DIPB, ENAL, ENAU, ENBL, ENBU, REGCEAL, REGCEAU, REGCEBL, REGCEBU, REGCLKAL, REGCLKAU, REGCLKBL, REGCLKBU, SSRAL, SSRAU, SSRBL, SSRBU, WEAL, WEAU, WEBL, WEBU) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [14:0] ADDRAU ;
input [14:0] ADDRBU ;
input [15:0] ADDRAL ;
input [15:0] ADDRBL ;
input CASCADEINLATA ;
input CASCADEINLATB ;
input CASCADEINREGA ;
input CASCADEINREGB ;
input CLKAL ;
input CLKAU ;
input CLKBL ;
input CLKBU ;
input [31:0] DIA ;
input [31:0] DIB ;
input [3:0] DIPA ;
input [3:0] DIPB ;
input ENAL ;
input ENAU ;
input ENBL ;
input ENBU ;
input REGCEAL ;
input REGCEAU ;
input REGCEBL ;
input REGCEBU ;
input REGCLKAL ;
input REGCLKAU ;
input REGCLKBL ;
input REGCLKBU ;
input SSRAL ;
input SSRAU ;
input SSRBL ;
input SSRBU ;
input [3:0] WEAL ;
input [3:0] WEAU ;
input [7:0] WEBL ;
input [7:0] WEBU ;
output CASCADEOUTLATA ;
output CASCADEOUTLATB ;
output CASCADEOUTREGA ;
output CASCADEOUTREGB ;
output [31:0] DOA ;
output [31:0] DOB ;
output [3:0] DOPA ;
output [3:0] DOPB ;
parameter DOA_REG = 0;
parameter DOB_REG = 0;
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_40 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_41 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_42 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_43 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_44 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_45 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_46 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_47 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_48 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_49 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_50 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_51 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_52 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_53 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_54 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_55 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_56 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_57 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_58 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_59 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_60 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_61 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_62 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_63 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_64 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_65 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_66 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_67 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_68 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_69 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_70 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_71 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_72 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_73 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_74 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_75 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_76 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_77 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_78 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_79 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 36'h0;
parameter INIT_B = 36'h0;
parameter INIT_FILE = "NONE";
parameter RAM_EXTENSION_A = "NONE";
parameter RAM_EXTENSION_B = "NONE";
parameter READ_WIDTH_A = 0;
parameter READ_WIDTH_B = 0;
parameter SIM_COLLISION_CHECK = "ALL";
parameter SIM_MODE = "SAFE";
parameter SRVAL_A = 36'h0;
parameter SRVAL_B = 36'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
parameter WRITE_WIDTH_A = 0;
parameter WRITE_WIDTH_B = 0;
endmodule
//#### END MODULE DEFINITION FOR: RAMB36_EXP ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S1 ###
module RAMB4_S1 (DO, ADDR, CLK, DI, EN, RST, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [11:0] ADDR ;
input [0:0] DI ;
input EN ;
input CLK ;
input WE ;
input RST ;
output [0:0] DO ;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S1 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S16 ###
module RAMB4_S16 (DO, ADDR, CLK, DI, EN, RST, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [7:0] ADDR ;
input [15:0] DI ;
input EN ;
input CLK ;
input WE ;
input RST ;
output [15:0] DO ;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S16 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S16_S16 ###
module RAMB4_S16_S16 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, RSTA, RSTB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [7:0] ADDRA ;
input [15:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input RSTA ;
input [7:0] ADDRB ;
input [15:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input RSTB ;
output [15:0] DOA ;
output [15:0] DOB ;
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S16_S16 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S1_S1 ###
module RAMB4_S1_S1 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, RSTA, RSTB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [11:0] ADDRA ;
input [0:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input RSTA ;
input [11:0] ADDRB ;
input [0:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input RSTB ;
output [0:0] DOA ;
output [0:0] DOB ;
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S1_S1 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S1_S16 ###
module RAMB4_S1_S16 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, RSTA, RSTB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [11:0] ADDRA ;
input [0:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input RSTA ;
input [7:0] ADDRB ;
input [15:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input RSTB ;
output [0:0] DOA ;
output [15:0] DOB ;
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S1_S16 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S1_S2 ###
module RAMB4_S1_S2 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, RSTA, RSTB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [11:0] ADDRA ;
input [0:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input RSTA ;
input [10:0] ADDRB ;
input [1:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input RSTB ;
output [0:0] DOA ;
output [1:0] DOB ;
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S1_S2 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S1_S4 ###
module RAMB4_S1_S4 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, RSTA, RSTB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [11:0] ADDRA ;
input [0:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input RSTA ;
input [9:0] ADDRB ;
input [3:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input RSTB ;
output [0:0] DOA ;
output [3:0] DOB ;
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S1_S4 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S1_S8 ###
module RAMB4_S1_S8 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, RSTA, RSTB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [11:0] ADDRA ;
input [0:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input RSTA ;
input [8:0] ADDRB ;
input [7:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input RSTB ;
output [0:0] DOA ;
output [7:0] DOB ;
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S1_S8 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S2 ###
module RAMB4_S2 (DO, ADDR, CLK, DI, EN, RST, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [10:0] ADDR ;
input [1:0] DI ;
input EN ;
input CLK ;
input WE ;
input RST ;
output [1:0] DO ;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S2 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S2_S16 ###
module RAMB4_S2_S16 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, RSTA, RSTB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [10:0] ADDRA ;
input [1:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input RSTA ;
input [7:0] ADDRB ;
input [15:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input RSTB ;
output [1:0] DOA ;
output [15:0] DOB ;
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S2_S16 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S2_S2 ###
module RAMB4_S2_S2 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, RSTA, RSTB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [10:0] ADDRA ;
input [1:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input RSTA ;
input [10:0] ADDRB ;
input [1:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input RSTB ;
output [1:0] DOA ;
output [1:0] DOB ;
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S2_S2 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S2_S4 ###
module RAMB4_S2_S4 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, RSTA, RSTB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [10:0] ADDRA ;
input [1:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input RSTA ;
input [9:0] ADDRB ;
input [3:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input RSTB ;
output [1:0] DOA ;
output [3:0] DOB ;
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S2_S4 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S2_S8 ###
module RAMB4_S2_S8 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, RSTA, RSTB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [10:0] ADDRA ;
input [1:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input RSTA ;
input [8:0] ADDRB ;
input [7:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input RSTB ;
output [1:0] DOA ;
output [7:0] DOB ;
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S2_S8 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S4 ###
module RAMB4_S4 (DO, ADDR, CLK, DI, EN, RST, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [9:0] ADDR ;
input [3:0] DI ;
input EN ;
input CLK ;
input WE ;
input RST ;
output [3:0] DO ;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S4 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S4_S16 ###
module RAMB4_S4_S16 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, RSTA, RSTB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [9:0] ADDRA ;
input [3:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input RSTA ;
input [7:0] ADDRB ;
input [15:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input RSTB ;
output [3:0] DOA ;
output [15:0] DOB ;
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S4_S16 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S4_S4 ###
module RAMB4_S4_S4 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, RSTA, RSTB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [9:0] ADDRA ;
input [3:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input RSTA ;
input [9:0] ADDRB ;
input [3:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input RSTB ;
output [3:0] DOA ;
output [3:0] DOB ;
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S4_S4 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S4_S8 ###
module RAMB4_S4_S8 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, RSTA, RSTB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [9:0] ADDRA ;
input [3:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input RSTA ;
input [8:0] ADDRB ;
input [7:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input RSTB ;
output [3:0] DOA ;
output [7:0] DOB ;
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S4_S8 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S8 ###
module RAMB4_S8 (DO, ADDR, CLK, DI, EN, RST, WE) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [8:0] ADDR ;
input [7:0] DI ;
input EN ;
input CLK ;
input WE ;
input RST ;
output [7:0] DO ;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S8 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S8_S16 ###
module RAMB4_S8_S16 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, RSTA, RSTB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [8:0] ADDRA ;
input [7:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input RSTA ;
input [7:0] ADDRB ;
input [15:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input RSTB ;
output [7:0] DOA ;
output [15:0] DOB ;
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S8_S16 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB4_S8_S8 ###
module RAMB4_S8_S8 (DOA, DOB, ADDRA, ADDRB, CLKA, CLKB, DIA, DIB, ENA, ENB, RSTA, RSTB, WEA, WEB) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [8:0] ADDRA ;
input [7:0] DIA ;
input ENA ;
input CLKA ;
input WEA ;
input RSTA ;
input [8:0] ADDRB ;
input [7:0] DIB ;
input ENB ;
input CLKB ;
input WEB ;
input RSTB ;
output [7:0] DOA ;
output [7:0] DOB ;
parameter SIM_COLLISION_CHECK = "ALL";
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: RAMB4_S8_S8 ####

//#### BEGIN MODULE DEFINITION FOR :RAMB8BWER ###
module RAMB8BWER (DOADO, DOBDO, DOPADOP, DOPBDOP, 
		  ADDRAWRADDR, ADDRBRDADDR, CLKAWRCLK, CLKBRDCLK, DIADI, DIBDI, DIPADIP, DIPBDIP, ENAWREN, ENBRDEN, REGCEA, REGCEBREGCE, RSTA, RSTBRST, WEAWEL, WEBWEU) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [12:0] ADDRAWRADDR ;
input [12:0] ADDRBRDADDR ;
input CLKAWRCLK ;
input CLKBRDCLK ;
input [15:0] DIADI ;
input [15:0] DIBDI ;
input [1:0] DIPADIP ;
input [1:0] DIPBDIP ;
input ENAWREN ;
input ENBRDEN ;
input REGCEA ;
input REGCEBREGCE ;
input RSTA ;
input RSTBRST ;
input [1:0] WEAWEL ;
input [1:0] WEBWEU ;
output [15:0] DOADO ;
output [15:0] DOBDO ;
output [1:0] DOPADOP ;
output [1:0] DOPBDOP ;
parameter DATA_WIDTH_A = 0;
parameter DATA_WIDTH_B = 0;
parameter DOA_REG = 0;
parameter DOB_REG = 0;
parameter EN_RSTRAM_A = "TRUE";
parameter EN_RSTRAM_B = "TRUE";
parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 18'h0;
parameter INIT_B = 18'h0;
parameter INIT_FILE = "NONE";
parameter RAM_MODE = "TDP";
parameter RSTTYPE = "SYNC";
parameter RST_PRIORITY_A = "CE";
parameter RST_PRIORITY_B = "CE";
parameter SETUP_ALL = 1000;
parameter SETUP_READ_FIRST = 3000;
parameter SIM_COLLISION_CHECK = "ALL";
parameter SRVAL_A = 18'h0;
parameter SRVAL_B = 18'h0;
parameter WRITE_MODE_A = "WRITE_FIRST";
parameter WRITE_MODE_B = "WRITE_FIRST";
endmodule
//#### END MODULE DEFINITION FOR: RAMB8BWER ####

//#### BEGIN MODULE DEFINITION FOR :ROM128X1 ###
module ROM128X1 (O, A0, A1, A2, A3, A4, A5, A6) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input A5 ;
input A6 ;
output O ;
parameter INIT = 128'h00000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: ROM128X1 ####

//#### BEGIN MODULE DEFINITION FOR :ROM16X1 ###
module ROM16X1 (O, A0, A1, A2, A3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
output O ;
parameter INIT = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: ROM16X1 ####

//#### BEGIN MODULE DEFINITION FOR :ROM256X1 ###
module ROM256X1 (O, A0, A1, A2, A3, A4, A5, A6, A7) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input A5 ;
input A6 ;
input A7 ;
output O ;
parameter INIT = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: ROM256X1 ####

//#### BEGIN MODULE DEFINITION FOR :ROM32X1 ###
module ROM32X1 (O, A0, A1, A2, A3, A4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
output O ;
parameter INIT = 32'h00000000;
endmodule
//#### END MODULE DEFINITION FOR: ROM32X1 ####

//#### BEGIN MODULE DEFINITION FOR :ROM64X1 ###
module ROM64X1 (O, A0, A1, A2, A3, A4, A5) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input A4 ;
input A5 ;
output O ;
parameter INIT = 64'h0000000000000000;
endmodule
//#### END MODULE DEFINITION FOR: ROM64X1 ####

//#### BEGIN MODULE DEFINITION FOR :SIM_CONFIGE2 ###
module SIM_CONFIGE2 ( 
                   CSOB,
                   DONE,
                   CCLK,
                   CSB,
                   D,
                   INITB,
                   M,
                   PROGB,
                   RDWRB
                   ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CCLK ;
input CSB ;
input [2:0] M ;
input PROGB ;
input RDWRB ;
output CSOB ;
inout DONE ;
inout [31:0] D ;
inout INITB ;
parameter DEVICE_ID = 32'h0;
parameter ICAP_SUPPORT = "FALSE";
parameter ICAP_WIDTH = "X8";
endmodule
//#### END MODULE DEFINITION FOR: SIM_CONFIGE2 ####

//#### BEGIN MODULE DEFINITION FOR :SIM_CONFIG_S3A ###
module SIM_CONFIG_S3A (
                   CSOB,
                   DONE,
                   CCLK,
                   D,
                   DCMLOCK,
                   CSIB,
                   INITB,
                   M,
                   PROGB,
                   RDWRB
                   ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CCLK ;
input DCMLOCK ;
input CSIB ;
input [2:0] M ;
input PROGB ;
input RDWRB ;
output CSOB ;
inout DONE ;
inout [7:0] D ;
inout INITB ;
parameter DEVICE_ID = 32'h0;
endmodule
//#### END MODULE DEFINITION FOR: SIM_CONFIG_S3A ####

//#### BEGIN MODULE DEFINITION FOR :SIM_CONFIG_S3A_SERIAL ###
module SIM_CONFIG_S3A_SERIAL (
                   DONE,
                   CCLK,
                   DIN,
                   INITB,
                   M,
                   PROGB
                   ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CCLK ;
input DIN ;
input [2:0] M ;
input PROGB ;
inout DONE ;
inout INITB ;
parameter DEVICE_ID = 32'h0;
endmodule
//#### END MODULE DEFINITION FOR: SIM_CONFIG_S3A_SERIAL ####

//#### BEGIN MODULE DEFINITION FOR :SIM_CONFIG_S6 ###
module SIM_CONFIG_S6 (
                   BUSY,
                   CSOB,
                   DONE,
                   CCLK,
                   D,
                   CSIB,
                   INITB,
                   M,
                   PROGB,
                   RDWRB
                   ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CCLK ;
input CSIB ;
input [1:0] M ;
input PROGB ;
input RDWRB ;
output BUSY ;
output CSOB ;
inout DONE ;
inout [15:0] D ;
inout INITB ;
parameter cfg_Tprog = 500000;
parameter cfg_Tpl = 5000000;
parameter DEVICE_ID = 32'h0;
parameter ICAP_SUPPORT = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: SIM_CONFIG_S6 ####

//#### BEGIN MODULE DEFINITION FOR :SIM_CONFIG_S6_SERIAL ###
module SIM_CONFIG_S6_SERIAL (
                   DONE,
                   CCLK,
                   DIN,
                   INITB,
                   M,
                   PROGB
                   ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CCLK ;
input DIN ;
input [1:0] M ;
input PROGB ;
inout DONE ;
inout INITB ;
parameter DEVICE_ID = 32'h0;
endmodule
//#### END MODULE DEFINITION FOR: SIM_CONFIG_S6_SERIAL ####

//#### BEGIN MODULE DEFINITION FOR :SIM_CONFIG_V5 ###
module SIM_CONFIG_V5 ( BUSY,
                   CSOB,
                   DONE,
                   CCLK,
                   CSB,
                   D,
                   DCMLOCK,
                   INITB,
                   M,
                   PROGB,
                   RDWRB
                   ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CCLK ;
input CSB ;
input DCMLOCK ;
input [2:0] M ;
input PROGB ;
input RDWRB ;
output BUSY ;
output CSOB ;
inout DONE ;
inout [31:0] D ;
inout INITB ;
parameter DEVICE_ID = 32'h0;
endmodule
//#### END MODULE DEFINITION FOR: SIM_CONFIG_V5 ####

//#### BEGIN MODULE DEFINITION FOR :SIM_CONFIG_V5_SERIAL ###
module SIM_CONFIG_V5_SERIAL (
                   DONE,
                   DOUT,
                   CCLK,
                   DIN,
                   INITB,
                   M,
                   PROGB
                   ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CCLK ;
input DIN ;
input [2:0] M ;
input PROGB ;
output DOUT ;
inout DONE ;
inout INITB ;
parameter DEVICE_ID = 32'h0;
endmodule
//#### END MODULE DEFINITION FOR: SIM_CONFIG_V5_SERIAL ####

//#### BEGIN MODULE DEFINITION FOR :SIM_CONFIG_V6 ###
module SIM_CONFIG_V6 ( BUSY,
                   CSOB,
                   DONE,
                   CCLK,
                   CSB,
                   D,
                   INITB,
                   M,
                   PROGB,
                   RDWRB
                   ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CCLK ;
input CSB ;
input [2:0] M ;
input PROGB ;
input RDWRB ;
output BUSY ;
output CSOB ;
inout DONE ;
inout [31:0] D ;
inout INITB ;
parameter DEVICE_ID = 32'h0;
parameter ICAP_SUPPORT = "FALSE";
parameter ICAP_WIDTH = "X8";
endmodule
//#### END MODULE DEFINITION FOR: SIM_CONFIG_V6 ####

//#### BEGIN MODULE DEFINITION FOR :SIM_CONFIG_V6_SERIAL ###
module SIM_CONFIG_V6_SERIAL ( 
                   DONE,
                   DOUT,
                   CCLK,
                   DIN,
                   INITB,
                   M,
                   PROGB
                   ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CCLK ;
input DIN ;
input [2:0] M ;
input PROGB ;
output DOUT ;
inout DONE ;
inout INITB ;
parameter DEVICE_ID = 32'h0;
endmodule
//#### END MODULE DEFINITION FOR: SIM_CONFIG_V6_SERIAL ####

//#### BEGIN MODULE DEFINITION FOR :SPI_ACCESS ###
module SPI_ACCESS (
   MISO,
   CLK,
   CSB,
   MOSI
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLK ;
input CSB ;
input MOSI ;
output MISO ;
parameter SIM_DELAY_TYPE = "SCALED";
parameter SIM_DEVICE = "3S1400AN";
parameter SIM_FACTORY_ID = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
parameter SIM_USER_ID =    512'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
parameter SIM_MEM_FILE = "NONE";
endmodule
//#### END MODULE DEFINITION FOR: SPI_ACCESS ####

//#### BEGIN MODULE DEFINITION FOR :SRL16 ###
module SRL16 (Q, A0, A1, A2, A3, CLK, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input CLK ;
input D ;
output Q ;
parameter INIT = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: SRL16 ####

//#### BEGIN MODULE DEFINITION FOR :SRL16E ###
module SRL16E (Q, A0, A1, A2, A3, CE, CLK, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input CE ;
input CLK ;
input D ;
output Q ;
parameter INIT = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: SRL16E ####

//#### BEGIN MODULE DEFINITION FOR :SRL16E_1 ###
module SRL16E_1 (Q, A0, A1, A2, A3, CE, CLK, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input CE ;
input CLK ;
input D ;
output Q ;
parameter INIT = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: SRL16E_1 ####

//#### BEGIN MODULE DEFINITION FOR :SRL16_1 ###
module SRL16_1 (Q, A0, A1, A2, A3, CLK, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input CLK ;
input D ;
output Q ;
parameter INIT = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: SRL16_1 ####

//#### BEGIN MODULE DEFINITION FOR :SRLC16 ###
module SRLC16 (Q, Q15, A0, A1, A2, A3, CLK, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input CLK ;
input D ;
output Q ;
output Q15 ;
parameter INIT = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: SRLC16 ####

//#### BEGIN MODULE DEFINITION FOR :SRLC16E ###
module SRLC16E (Q, Q15, A0, A1, A2, A3, CE, CLK, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input CE ;
input CLK ;
input D ;
output Q ;
output Q15 ;
parameter INIT = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: SRLC16E ####

//#### BEGIN MODULE DEFINITION FOR :SRLC16E_1 ###
module SRLC16E_1 (Q, Q15, A0, A1, A2, A3, CE, CLK, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input CE ;
input CLK ;
input D ;
output Q ;
output Q15 ;
parameter INIT = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: SRLC16E_1 ####

//#### BEGIN MODULE DEFINITION FOR :SRLC16_1 ###
module SRLC16_1 (Q, Q15, A0, A1, A2, A3, CLK, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input A0 ;
input A1 ;
input A2 ;
input A3 ;
input CLK ;
input D ;
output Q ;
output Q15 ;
parameter INIT = 16'h0000;
endmodule
//#### END MODULE DEFINITION FOR: SRLC16_1 ####

//#### BEGIN MODULE DEFINITION FOR :SRLC32E ###
module SRLC32E (Q, Q31, A, CE, CLK, D) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input [4:0] A ;
input CE ;
input CLK ;
input D ;
output Q ;
output Q31 ;
parameter INIT = 32'h00000000;
endmodule
//#### END MODULE DEFINITION FOR: SRLC32E ####

//#### BEGIN MODULE DEFINITION FOR :STARTUPE2 ###
module STARTUPE2 (
  CFGCLK,
  CFGMCLK,
  EOS,
  PREQ,

  CLK,
  GSR,
  GTS,
  KEYCLEARB,
  PACK,
  USRCCLKO,
  USRCCLKTS,
  USRDONEO,
  USRDONETS
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLK ;
input GSR ;
input GTS ;
input KEYCLEARB ;
input PACK ;
input USRCCLKO ;
input USRCCLKTS ;
input USRDONEO ;
input USRDONETS ;
output CFGCLK ;
output CFGMCLK ;
output EOS ;
output PREQ ;
parameter PROG_USR = "FALSE";
parameter SIM_CCLK_FREQ = 0.0;
endmodule
//#### END MODULE DEFINITION FOR: STARTUPE2 ####

//#### BEGIN MODULE DEFINITION FOR :STARTUP_FPGACORE ###
module STARTUP_FPGACORE (CLK, GSR) /* synthesis syn_black_box  syn_lib_cell=1
 .noprune=1
 */;
input CLK ;
input GSR ;
endmodule
//#### END MODULE DEFINITION FOR: STARTUP_FPGACORE ####

//#### BEGIN MODULE DEFINITION FOR :STARTUP_SPARTAN3 ###
module STARTUP_SPARTAN3 (CLK, GSR, GTS) /* synthesis syn_black_box  syn_lib_cell=1
 .noprune=1
 */;
input CLK ;
input GSR ;
input GTS ;
endmodule
//#### END MODULE DEFINITION FOR: STARTUP_SPARTAN3 ####

//#### BEGIN MODULE DEFINITION FOR :STARTUP_SPARTAN3A ###
module STARTUP_SPARTAN3A (CLK, GSR, GTS) /* synthesis syn_black_box  syn_lib_cell=1
 .noprune=1
 */;
input CLK ;
input GSR ;
input GTS ;
endmodule
//#### END MODULE DEFINITION FOR: STARTUP_SPARTAN3A ####

//#### BEGIN MODULE DEFINITION FOR :STARTUP_SPARTAN3E ###
module STARTUP_SPARTAN3E (CLK, GSR, GTS, MBT) /* synthesis syn_black_box  syn_lib_cell=1
 .noprune=1
 */;
input CLK ;
input GSR ;
input GTS ;
input MBT ;
endmodule
//#### END MODULE DEFINITION FOR: STARTUP_SPARTAN3E ####

//#### BEGIN MODULE DEFINITION FOR :STARTUP_SPARTAN6 ###
module STARTUP_SPARTAN6 (
  CFGCLK,
  CFGMCLK,
  EOS,
  CLK,
  GSR,
  GTS,
  KEYCLEARB
) /* synthesis syn_black_box  syn_lib_cell=1
 .noprune=1
 */;
input CLK ;
input GSR ;
input GTS ;
input KEYCLEARB ;
output CFGCLK ;
output CFGMCLK ;
output EOS ;
endmodule
//#### END MODULE DEFINITION FOR: STARTUP_SPARTAN6 ####

//#### BEGIN MODULE DEFINITION FOR :STARTUP_VIRTEX4 ###
module STARTUP_VIRTEX4 (EOS, CLK, GSR, GTS, USRCCLKO, USRCCLKTS, USRDONEO, USRDONETS) /* synthesis syn_black_box  syn_lib_cell=1
 .noprune=1
 */;
input CLK ;
input GSR ;
input GTS ;
input USRCCLKO ;
input USRCCLKTS ;
input USRDONEO ;
input USRDONETS ;
output EOS ;
endmodule
//#### END MODULE DEFINITION FOR: STARTUP_VIRTEX4 ####

//#### BEGIN MODULE DEFINITION FOR :STARTUP_VIRTEX5 ###
module STARTUP_VIRTEX5 (
        CFGCLK,
        CFGMCLK,
        DINSPI,
	EOS,
        TCKSPI,
	CLK,
	GSR,
	GTS,
	USRCCLKO,
	USRCCLKTS,
	USRDONEO,
	USRDONETS
) /* synthesis syn_black_box  syn_lib_cell=1
 .noprune=1
 */;
input CLK ;
input GSR ;
input GTS ;
input USRCCLKO ;
input USRCCLKTS ;
input USRDONEO ;
input USRDONETS ;
output CFGCLK ;
output CFGMCLK ;
output DINSPI ;
output EOS ;
output TCKSPI ;
endmodule
//#### END MODULE DEFINITION FOR: STARTUP_VIRTEX5 ####

//#### BEGIN MODULE DEFINITION FOR :STARTUP_VIRTEX6 ###
module STARTUP_VIRTEX6 (
  CFGCLK,
  CFGMCLK,
  DINSPI,
  EOS,
  PREQ,
  TCKSPI,
  CLK,
  GSR,
  GTS,
  KEYCLEARB,
  PACK,
  USRCCLKO,
  USRCCLKTS,
  USRDONEO,
  USRDONETS
) /* synthesis syn_black_box  syn_lib_cell=1
 .noprune=1
 */;
input CLK ;
input GSR ;
input GTS ;
input KEYCLEARB ;
input PACK ;
input USRCCLKO ;
input USRCCLKTS ;
input USRDONEO ;
input USRDONETS ;
output CFGCLK ;
output CFGMCLK ;
output DINSPI ;
output EOS ;
output PREQ ;
output TCKSPI ;
parameter PROG_USR = "FALSE";
endmodule
//#### END MODULE DEFINITION FOR: STARTUP_VIRTEX6 ####

//#### BEGIN MODULE DEFINITION FOR :SUSPEND_SYNC ###
module SUSPEND_SYNC (
  SREQ,
  CLK,
  SACK
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLK ;
input SACK ;
output SREQ ;
endmodule
//#### END MODULE DEFINITION FOR: SUSPEND_SYNC ####

//#### BEGIN MODULE DEFINITION FOR :SYSMON ###
module SYSMON (
        ALM,
        BUSY,
        CHANNEL,
        DO,
        DRDY,
        EOC,
        EOS,
        JTAGBUSY,
        JTAGLOCKED,
        JTAGMODIFIED,
        OT,
        CONVST,
        CONVSTCLK,
        DADDR,
        DCLK,
        DEN,
        DI,
        DWE,
        RESET,
        VAUXN,
        VAUXP,
        VN,
        VP

) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CONVST ;
input CONVSTCLK ;
input DCLK ;
input DEN ;
input DWE ;
input RESET ;
input VN ;
input VP ;
input [15:0] DI ;
input [15:0] VAUXN ;
input [15:0] VAUXP ;
input [6:0] DADDR ;
output BUSY ;
output DRDY ;
output EOC ;
output EOS ;
output JTAGBUSY ;
output JTAGLOCKED ;
output JTAGMODIFIED ;
output OT ;
output [15:0] DO ;
output [2:0] ALM ;
output [4:0] CHANNEL ;
parameter  [15:0] INIT_40 = 16'h0;
parameter  [15:0] INIT_41 = 16'h0;
parameter  [15:0] INIT_42 = 16'h0800;
parameter  [15:0] INIT_43 = 16'h0;
parameter  [15:0] INIT_44 = 16'h0;
parameter  [15:0] INIT_45 = 16'h0;
parameter  [15:0] INIT_46 = 16'h0;
parameter  [15:0] INIT_47 = 16'h0;
parameter  [15:0] INIT_48 = 16'h0;
parameter  [15:0] INIT_49 = 16'h0;
parameter  [15:0] INIT_4A = 16'h0;
parameter  [15:0] INIT_4B = 16'h0;
parameter  [15:0] INIT_4C = 16'h0;
parameter  [15:0] INIT_4D = 16'h0;
parameter  [15:0] INIT_4E = 16'h0;
parameter  [15:0] INIT_4F = 16'h0;
parameter  [15:0] INIT_50 = 16'h0;
parameter  [15:0] INIT_51 = 16'h0;
parameter  [15:0] INIT_52 = 16'h0;
parameter  [15:0] INIT_53 = 16'h0;
parameter  [15:0] INIT_54 = 16'h0;
parameter  [15:0] INIT_55 = 16'h0;
parameter  [15:0] INIT_56 = 16'h0;
parameter  [15:0] INIT_57 = 16'h0;
parameter SIM_DEVICE = "VIRTEX5";
parameter SIM_MONITOR_FILE = "design.txt";
endmodule
//#### END MODULE DEFINITION FOR: SYSMON ####

//#### BEGIN MODULE DEFINITION FOR :TBLOCK ###
module TBLOCK () /* synthesis syn_black_box  syn_lib_cell=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: TBLOCK ####

//#### BEGIN MODULE DEFINITION FOR :TEMAC ###
module TEMAC (
	DCRHOSTDONEIR,
	EMAC0CLIENTANINTERRUPT,
	EMAC0CLIENTRXBADFRAME,
	EMAC0CLIENTRXCLIENTCLKOUT,
	EMAC0CLIENTRXD,
	EMAC0CLIENTRXDVLD,
	EMAC0CLIENTRXDVLDMSW,
	EMAC0CLIENTRXFRAMEDROP,
	EMAC0CLIENTRXGOODFRAME,
	EMAC0CLIENTRXSTATS,
	EMAC0CLIENTRXSTATSBYTEVLD,
	EMAC0CLIENTRXSTATSVLD,
	EMAC0CLIENTTXACK,
	EMAC0CLIENTTXCLIENTCLKOUT,
	EMAC0CLIENTTXCOLLISION,
	EMAC0CLIENTTXRETRANSMIT,
	EMAC0CLIENTTXSTATS,
	EMAC0CLIENTTXSTATSBYTEVLD,
	EMAC0CLIENTTXSTATSVLD,
	EMAC0PHYENCOMMAALIGN,
	EMAC0PHYLOOPBACKMSB,
	EMAC0PHYMCLKOUT,
	EMAC0PHYMDOUT,
	EMAC0PHYMDTRI,
	EMAC0PHYMGTRXRESET,
	EMAC0PHYMGTTXRESET,
	EMAC0PHYPOWERDOWN,
	EMAC0PHYSYNCACQSTATUS,
	EMAC0PHYTXCHARDISPMODE,
	EMAC0PHYTXCHARDISPVAL,
	EMAC0PHYTXCHARISK,
	EMAC0PHYTXCLK,
	EMAC0PHYTXD,
	EMAC0PHYTXEN,
	EMAC0PHYTXER,
	EMAC0PHYTXGMIIMIICLKOUT,
	EMAC0SPEEDIS10100,
	EMAC1CLIENTANINTERRUPT,
	EMAC1CLIENTRXBADFRAME,
	EMAC1CLIENTRXCLIENTCLKOUT,
	EMAC1CLIENTRXD,
	EMAC1CLIENTRXDVLD,
	EMAC1CLIENTRXDVLDMSW,
	EMAC1CLIENTRXFRAMEDROP,
	EMAC1CLIENTRXGOODFRAME,
	EMAC1CLIENTRXSTATS,
	EMAC1CLIENTRXSTATSBYTEVLD,
	EMAC1CLIENTRXSTATSVLD,
	EMAC1CLIENTTXACK,
	EMAC1CLIENTTXCLIENTCLKOUT,
	EMAC1CLIENTTXCOLLISION,
	EMAC1CLIENTTXRETRANSMIT,
	EMAC1CLIENTTXSTATS,
	EMAC1CLIENTTXSTATSBYTEVLD,
	EMAC1CLIENTTXSTATSVLD,
	EMAC1PHYENCOMMAALIGN,
	EMAC1PHYLOOPBACKMSB,
	EMAC1PHYMCLKOUT,
	EMAC1PHYMDOUT,
	EMAC1PHYMDTRI,
	EMAC1PHYMGTRXRESET,
	EMAC1PHYMGTTXRESET,
	EMAC1PHYPOWERDOWN,
	EMAC1PHYSYNCACQSTATUS,
	EMAC1PHYTXCHARDISPMODE,
	EMAC1PHYTXCHARDISPVAL,
	EMAC1PHYTXCHARISK,
	EMAC1PHYTXCLK,
	EMAC1PHYTXD,
	EMAC1PHYTXEN,
	EMAC1PHYTXER,
	EMAC1PHYTXGMIIMIICLKOUT,
	EMAC1SPEEDIS10100,
	EMACDCRACK,
	EMACDCRDBUS,
	HOSTMIIMRDY,
	HOSTRDDATA,

	CLIENTEMAC0DCMLOCKED,
	CLIENTEMAC0PAUSEREQ,
	CLIENTEMAC0PAUSEVAL,
	CLIENTEMAC0RXCLIENTCLKIN,
	CLIENTEMAC0TXCLIENTCLKIN,
	CLIENTEMAC0TXD,
	CLIENTEMAC0TXDVLD,
	CLIENTEMAC0TXDVLDMSW,
	CLIENTEMAC0TXFIRSTBYTE,
	CLIENTEMAC0TXIFGDELAY,
	CLIENTEMAC0TXUNDERRUN,
	CLIENTEMAC1DCMLOCKED,
	CLIENTEMAC1PAUSEREQ,
	CLIENTEMAC1PAUSEVAL,
	CLIENTEMAC1RXCLIENTCLKIN,
	CLIENTEMAC1TXCLIENTCLKIN,
	CLIENTEMAC1TXD,
	CLIENTEMAC1TXDVLD,
	CLIENTEMAC1TXDVLDMSW,
	CLIENTEMAC1TXFIRSTBYTE,
	CLIENTEMAC1TXIFGDELAY,
	CLIENTEMAC1TXUNDERRUN,
	DCREMACABUS,
	DCREMACCLK,
	DCREMACDBUS,
	DCREMACENABLE,
	DCREMACREAD,
	DCREMACWRITE,
	HOSTADDR,
	HOSTCLK,
	HOSTEMAC1SEL,
	HOSTMIIMSEL,
	HOSTOPCODE,
	HOSTREQ,
	HOSTWRDATA,
	PHYEMAC0COL,
	PHYEMAC0CRS,
	PHYEMAC0GTXCLK,
	PHYEMAC0MCLKIN,
	PHYEMAC0MDIN,
	PHYEMAC0MIITXCLK,
	PHYEMAC0PHYAD,
	PHYEMAC0RXBUFERR,
	PHYEMAC0RXBUFSTATUS,
	PHYEMAC0RXCHARISCOMMA,
	PHYEMAC0RXCHARISK,
	PHYEMAC0RXCHECKINGCRC,
	PHYEMAC0RXCLK,
	PHYEMAC0RXCLKCORCNT,
	PHYEMAC0RXCOMMADET,
	PHYEMAC0RXD,
	PHYEMAC0RXDISPERR,
	PHYEMAC0RXDV,
	PHYEMAC0RXER,
	PHYEMAC0RXLOSSOFSYNC,
	PHYEMAC0RXNOTINTABLE,
	PHYEMAC0RXRUNDISP,
	PHYEMAC0SIGNALDET,
	PHYEMAC0TXBUFERR,
	PHYEMAC0TXGMIIMIICLKIN,
	PHYEMAC1COL,
	PHYEMAC1CRS,
	PHYEMAC1GTXCLK,
	PHYEMAC1MCLKIN,
	PHYEMAC1MDIN,
	PHYEMAC1MIITXCLK,
	PHYEMAC1PHYAD,
	PHYEMAC1RXBUFERR,
	PHYEMAC1RXBUFSTATUS,
	PHYEMAC1RXCHARISCOMMA,
	PHYEMAC1RXCHARISK,
	PHYEMAC1RXCHECKINGCRC,
	PHYEMAC1RXCLK,
	PHYEMAC1RXCLKCORCNT,
	PHYEMAC1RXCOMMADET,
	PHYEMAC1RXD,
	PHYEMAC1RXDISPERR,
	PHYEMAC1RXDV,
	PHYEMAC1RXER,
	PHYEMAC1RXLOSSOFSYNC,
	PHYEMAC1RXNOTINTABLE,
	PHYEMAC1RXRUNDISP,
	PHYEMAC1SIGNALDET,
	PHYEMAC1TXBUFERR,
	PHYEMAC1TXGMIIMIICLKIN,
	RESET

) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLIENTEMAC0DCMLOCKED ;
input CLIENTEMAC0PAUSEREQ ;
input CLIENTEMAC0RXCLIENTCLKIN ;
input CLIENTEMAC0TXCLIENTCLKIN ;
input CLIENTEMAC0TXDVLD ;
input CLIENTEMAC0TXDVLDMSW ;
input CLIENTEMAC0TXFIRSTBYTE ;
input CLIENTEMAC0TXUNDERRUN ;
input CLIENTEMAC1DCMLOCKED ;
input CLIENTEMAC1PAUSEREQ ;
input CLIENTEMAC1RXCLIENTCLKIN ;
input CLIENTEMAC1TXCLIENTCLKIN ;
input CLIENTEMAC1TXDVLD ;
input CLIENTEMAC1TXDVLDMSW ;
input CLIENTEMAC1TXFIRSTBYTE ;
input CLIENTEMAC1TXUNDERRUN ;
input DCREMACCLK ;
input DCREMACENABLE ;
input DCREMACREAD ;
input DCREMACWRITE ;
input HOSTCLK ;
input HOSTEMAC1SEL ;
input HOSTMIIMSEL ;
input HOSTREQ ;
input PHYEMAC0COL ;
input PHYEMAC0CRS ;
input PHYEMAC0GTXCLK ;
input PHYEMAC0MCLKIN ;
input PHYEMAC0MDIN ;
input PHYEMAC0MIITXCLK ;
input PHYEMAC0RXBUFERR ;
input PHYEMAC0RXCHARISCOMMA ;
input PHYEMAC0RXCHARISK ;
input PHYEMAC0RXCHECKINGCRC ;
input PHYEMAC0RXCLK ;
input PHYEMAC0RXCOMMADET ;
input PHYEMAC0RXDISPERR ;
input PHYEMAC0RXDV ;
input PHYEMAC0RXER ;
input PHYEMAC0RXNOTINTABLE ;
input PHYEMAC0RXRUNDISP ;
input PHYEMAC0SIGNALDET ;
input PHYEMAC0TXBUFERR ;
input PHYEMAC0TXGMIIMIICLKIN ;
input PHYEMAC1COL ;
input PHYEMAC1CRS ;
input PHYEMAC1GTXCLK ;
input PHYEMAC1MCLKIN ;
input PHYEMAC1MDIN ;
input PHYEMAC1MIITXCLK ;
input PHYEMAC1RXBUFERR ;
input PHYEMAC1RXCHARISCOMMA ;
input PHYEMAC1RXCHARISK ;
input PHYEMAC1RXCHECKINGCRC ;
input PHYEMAC1RXCLK ;
input PHYEMAC1RXCOMMADET ;
input PHYEMAC1RXDISPERR ;
input PHYEMAC1RXDV ;
input PHYEMAC1RXER ;
input PHYEMAC1RXNOTINTABLE ;
input PHYEMAC1RXRUNDISP ;
input PHYEMAC1SIGNALDET ;
input PHYEMAC1TXBUFERR ;
input PHYEMAC1TXGMIIMIICLKIN ;
input RESET ;
input [0:31] DCREMACDBUS ;
input [0:9] DCREMACABUS ;
input [15:0] CLIENTEMAC0PAUSEVAL ;
input [15:0] CLIENTEMAC0TXD ;
input [15:0] CLIENTEMAC1PAUSEVAL ;
input [15:0] CLIENTEMAC1TXD ;
input [1:0] HOSTOPCODE ;
input [1:0] PHYEMAC0RXBUFSTATUS ;
input [1:0] PHYEMAC0RXLOSSOFSYNC ;
input [1:0] PHYEMAC1RXBUFSTATUS ;
input [1:0] PHYEMAC1RXLOSSOFSYNC ;
input [2:0] PHYEMAC0RXCLKCORCNT ;
input [2:0] PHYEMAC1RXCLKCORCNT ;
input [31:0] HOSTWRDATA ;
input [4:0] PHYEMAC0PHYAD ;
input [4:0] PHYEMAC1PHYAD ;
input [7:0] CLIENTEMAC0TXIFGDELAY ;
input [7:0] CLIENTEMAC1TXIFGDELAY ;
input [7:0] PHYEMAC0RXD ;
input [7:0] PHYEMAC1RXD ;
input [9:0] HOSTADDR ;
output DCRHOSTDONEIR ;
output EMAC0CLIENTANINTERRUPT ;
output EMAC0CLIENTRXBADFRAME ;
output EMAC0CLIENTRXCLIENTCLKOUT ;
output EMAC0CLIENTRXDVLD ;
output EMAC0CLIENTRXDVLDMSW ;
output EMAC0CLIENTRXFRAMEDROP ;
output EMAC0CLIENTRXGOODFRAME ;
output EMAC0CLIENTRXSTATSBYTEVLD ;
output EMAC0CLIENTRXSTATSVLD ;
output EMAC0CLIENTTXACK ;
output EMAC0CLIENTTXCLIENTCLKOUT ;
output EMAC0CLIENTTXCOLLISION ;
output EMAC0CLIENTTXRETRANSMIT ;
output EMAC0CLIENTTXSTATS ;
output EMAC0CLIENTTXSTATSBYTEVLD ;
output EMAC0CLIENTTXSTATSVLD ;
output EMAC0PHYENCOMMAALIGN ;
output EMAC0PHYLOOPBACKMSB ;
output EMAC0PHYMCLKOUT ;
output EMAC0PHYMDOUT ;
output EMAC0PHYMDTRI ;
output EMAC0PHYMGTRXRESET ;
output EMAC0PHYMGTTXRESET ;
output EMAC0PHYPOWERDOWN ;
output EMAC0PHYSYNCACQSTATUS ;
output EMAC0PHYTXCHARDISPMODE ;
output EMAC0PHYTXCHARDISPVAL ;
output EMAC0PHYTXCHARISK ;
output EMAC0PHYTXCLK ;
output EMAC0PHYTXEN ;
output EMAC0PHYTXER ;
output EMAC0PHYTXGMIIMIICLKOUT ;
output EMAC0SPEEDIS10100 ;
output EMAC1CLIENTANINTERRUPT ;
output EMAC1CLIENTRXBADFRAME ;
output EMAC1CLIENTRXCLIENTCLKOUT ;
output EMAC1CLIENTRXDVLD ;
output EMAC1CLIENTRXDVLDMSW ;
output EMAC1CLIENTRXFRAMEDROP ;
output EMAC1CLIENTRXGOODFRAME ;
output EMAC1CLIENTRXSTATSBYTEVLD ;
output EMAC1CLIENTRXSTATSVLD ;
output EMAC1CLIENTTXACK ;
output EMAC1CLIENTTXCLIENTCLKOUT ;
output EMAC1CLIENTTXCOLLISION ;
output EMAC1CLIENTTXRETRANSMIT ;
output EMAC1CLIENTTXSTATS ;
output EMAC1CLIENTTXSTATSBYTEVLD ;
output EMAC1CLIENTTXSTATSVLD ;
output EMAC1PHYENCOMMAALIGN ;
output EMAC1PHYLOOPBACKMSB ;
output EMAC1PHYMCLKOUT ;
output EMAC1PHYMDOUT ;
output EMAC1PHYMDTRI ;
output EMAC1PHYMGTRXRESET ;
output EMAC1PHYMGTTXRESET ;
output EMAC1PHYPOWERDOWN ;
output EMAC1PHYSYNCACQSTATUS ;
output EMAC1PHYTXCHARDISPMODE ;
output EMAC1PHYTXCHARDISPVAL ;
output EMAC1PHYTXCHARISK ;
output EMAC1PHYTXCLK ;
output EMAC1PHYTXEN ;
output EMAC1PHYTXER ;
output EMAC1PHYTXGMIIMIICLKOUT ;
output EMAC1SPEEDIS10100 ;
output EMACDCRACK ;
output HOSTMIIMRDY ;
output [0:31] EMACDCRDBUS ;
output [15:0] EMAC0CLIENTRXD ;
output [15:0] EMAC1CLIENTRXD ;
output [31:0] HOSTRDDATA ;
output [6:0] EMAC0CLIENTRXSTATS ;
output [6:0] EMAC1CLIENTRXSTATS ;
output [7:0] EMAC0PHYTXD ;
output [7:0] EMAC1PHYTXD ;
parameter EMAC0_1000BASEX_ENABLE = "FALSE";
parameter EMAC0_ADDRFILTER_ENABLE = "FALSE";
parameter EMAC0_BYTEPHY = "FALSE";
parameter EMAC0_CONFIGVEC_79 = "FALSE";
parameter EMAC0_GTLOOPBACK = "FALSE";
parameter EMAC0_HOST_ENABLE = "FALSE";
parameter EMAC0_LTCHECK_DISABLE = "FALSE";
parameter EMAC0_MDIO_ENABLE = "FALSE";
parameter EMAC0_PHYINITAUTONEG_ENABLE = "FALSE";
parameter EMAC0_PHYISOLATE = "FALSE";
parameter EMAC0_PHYLOOPBACKMSB = "FALSE";
parameter EMAC0_PHYPOWERDOWN = "FALSE";
parameter EMAC0_PHYRESET = "FALSE";
parameter EMAC0_RGMII_ENABLE = "FALSE";
parameter EMAC0_RX16BITCLIENT_ENABLE = "FALSE";
parameter EMAC0_RXFLOWCTRL_ENABLE = "FALSE";
parameter EMAC0_RXHALFDUPLEX = "FALSE";
parameter EMAC0_RXINBANDFCS_ENABLE = "FALSE";
parameter EMAC0_RXJUMBOFRAME_ENABLE = "FALSE";
parameter EMAC0_RXRESET = "FALSE";
parameter EMAC0_RXVLAN_ENABLE = "FALSE";
parameter EMAC0_RX_ENABLE = "FALSE";
parameter EMAC0_SGMII_ENABLE = "FALSE";
parameter EMAC0_SPEED_LSB = "FALSE";
parameter EMAC0_SPEED_MSB = "FALSE";
parameter EMAC0_TX16BITCLIENT_ENABLE = "FALSE";
parameter EMAC0_TXFLOWCTRL_ENABLE = "FALSE";
parameter EMAC0_TXHALFDUPLEX = "FALSE";
parameter EMAC0_TXIFGADJUST_ENABLE = "FALSE";
parameter EMAC0_TXINBANDFCS_ENABLE = "FALSE";
parameter EMAC0_TXJUMBOFRAME_ENABLE = "FALSE";
parameter EMAC0_TXRESET = "FALSE";
parameter EMAC0_TXVLAN_ENABLE = "FALSE";
parameter EMAC0_TX_ENABLE = "FALSE";
parameter EMAC0_UNIDIRECTION_ENABLE = "FALSE";
parameter EMAC0_USECLKEN = "FALSE";
parameter EMAC1_1000BASEX_ENABLE = "FALSE";
parameter EMAC1_ADDRFILTER_ENABLE = "FALSE";
parameter EMAC1_BYTEPHY = "FALSE";
parameter EMAC1_CONFIGVEC_79 = "FALSE";
parameter EMAC1_GTLOOPBACK = "FALSE";
parameter EMAC1_HOST_ENABLE = "FALSE";
parameter EMAC1_LTCHECK_DISABLE = "FALSE";
parameter EMAC1_MDIO_ENABLE = "FALSE";
parameter EMAC1_PHYINITAUTONEG_ENABLE = "FALSE";
parameter EMAC1_PHYISOLATE = "FALSE";
parameter EMAC1_PHYLOOPBACKMSB = "FALSE";
parameter EMAC1_PHYPOWERDOWN = "FALSE";
parameter EMAC1_PHYRESET = "FALSE";
parameter EMAC1_RGMII_ENABLE = "FALSE";
parameter EMAC1_RX16BITCLIENT_ENABLE = "FALSE";
parameter EMAC1_RXFLOWCTRL_ENABLE = "FALSE";
parameter EMAC1_RXHALFDUPLEX = "FALSE";
parameter EMAC1_RXINBANDFCS_ENABLE = "FALSE";
parameter EMAC1_RXJUMBOFRAME_ENABLE = "FALSE";
parameter EMAC1_RXRESET = "FALSE";
parameter EMAC1_RXVLAN_ENABLE = "FALSE";
parameter EMAC1_RX_ENABLE = "FALSE";
parameter EMAC1_SGMII_ENABLE = "FALSE";
parameter EMAC1_SPEED_LSB = "FALSE";
parameter EMAC1_SPEED_MSB = "FALSE";
parameter EMAC1_TX16BITCLIENT_ENABLE = "FALSE";
parameter EMAC1_TXFLOWCTRL_ENABLE = "FALSE";
parameter EMAC1_TXHALFDUPLEX = "FALSE";
parameter EMAC1_TXIFGADJUST_ENABLE = "FALSE";
parameter EMAC1_TXINBANDFCS_ENABLE = "FALSE";
parameter EMAC1_TXJUMBOFRAME_ENABLE = "FALSE";
parameter EMAC1_TXRESET = "FALSE";
parameter EMAC1_TXVLAN_ENABLE = "FALSE";
parameter EMAC1_TX_ENABLE = "FALSE";
parameter EMAC1_UNIDIRECTION_ENABLE = "FALSE";
parameter EMAC1_USECLKEN = "FALSE";
parameter [0:7] EMAC0_DCRBASEADDR = 8'h00;
parameter [0:7] EMAC1_DCRBASEADDR = 8'h00;
parameter [47:0] EMAC0_PAUSEADDR = 48'h000000000000;
parameter [47:0] EMAC0_UNICASTADDR = 48'h000000000000;
parameter [47:0] EMAC1_PAUSEADDR = 48'h000000000000;
parameter [47:0] EMAC1_UNICASTADDR = 48'h000000000000;
parameter [8:0] EMAC0_LINKTIMERVAL = 9'h000;
parameter [8:0] EMAC1_LINKTIMERVAL = 9'h000;
endmodule
//#### END MODULE DEFINITION FOR: TEMAC ####

//#### BEGIN MODULE DEFINITION FOR :TEMAC_SINGLE ###
module TEMAC_SINGLE (
  DCRHOSTDONEIR,
  EMACCLIENTANINTERRUPT,
  EMACCLIENTRXBADFRAME,
  EMACCLIENTRXCLIENTCLKOUT,
  EMACCLIENTRXD,
  EMACCLIENTRXDVLD,
  EMACCLIENTRXDVLDMSW,
  EMACCLIENTRXFRAMEDROP,
  EMACCLIENTRXGOODFRAME,
  EMACCLIENTRXSTATS,
  EMACCLIENTRXSTATSBYTEVLD,
  EMACCLIENTRXSTATSVLD,
  EMACCLIENTTXACK,
  EMACCLIENTTXCLIENTCLKOUT,
  EMACCLIENTTXCOLLISION,
  EMACCLIENTTXRETRANSMIT,
  EMACCLIENTTXSTATS,
  EMACCLIENTTXSTATSBYTEVLD,
  EMACCLIENTTXSTATSVLD,
  EMACDCRACK,
  EMACDCRDBUS,
  EMACPHYENCOMMAALIGN,
  EMACPHYLOOPBACKMSB,
  EMACPHYMCLKOUT,
  EMACPHYMDOUT,
  EMACPHYMDTRI,
  EMACPHYMGTRXRESET,
  EMACPHYMGTTXRESET,
  EMACPHYPOWERDOWN,
  EMACPHYSYNCACQSTATUS,
  EMACPHYTXCHARDISPMODE,
  EMACPHYTXCHARDISPVAL,
  EMACPHYTXCHARISK,
  EMACPHYTXCLK,
  EMACPHYTXD,
  EMACPHYTXEN,
  EMACPHYTXER,
  EMACPHYTXGMIIMIICLKOUT,
  EMACSPEEDIS10100,
  HOSTMIIMRDY,
  HOSTRDDATA,
  CLIENTEMACDCMLOCKED,
  CLIENTEMACPAUSEREQ,
  CLIENTEMACPAUSEVAL,
  CLIENTEMACRXCLIENTCLKIN,
  CLIENTEMACTXCLIENTCLKIN,
  CLIENTEMACTXD,
  CLIENTEMACTXDVLD,
  CLIENTEMACTXDVLDMSW,
  CLIENTEMACTXFIRSTBYTE,
  CLIENTEMACTXIFGDELAY,
  CLIENTEMACTXUNDERRUN,
  DCREMACABUS,
  DCREMACCLK,
  DCREMACDBUS,
  DCREMACENABLE,
  DCREMACREAD,
  DCREMACWRITE,
  HOSTADDR,
  HOSTCLK,
  HOSTMIIMSEL,
  HOSTOPCODE,
  HOSTREQ,
  HOSTWRDATA,
  PHYEMACCOL,
  PHYEMACCRS,
  PHYEMACGTXCLK,
  PHYEMACMCLKIN,
  PHYEMACMDIN,
  PHYEMACMIITXCLK,
  PHYEMACPHYAD,
  PHYEMACRXBUFSTATUS,
  PHYEMACRXCHARISCOMMA,
  PHYEMACRXCHARISK,
  PHYEMACRXCLK,
  PHYEMACRXCLKCORCNT,
  PHYEMACRXD,
  PHYEMACRXDISPERR,
  PHYEMACRXDV,
  PHYEMACRXER,
  PHYEMACRXNOTINTABLE,
  PHYEMACRXRUNDISP,
  PHYEMACSIGNALDET,
  PHYEMACTXBUFERR,
  PHYEMACTXGMIIMIICLKIN,
  RESET
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CLIENTEMACDCMLOCKED ;
input CLIENTEMACPAUSEREQ ;
input CLIENTEMACRXCLIENTCLKIN ;
input CLIENTEMACTXCLIENTCLKIN ;
input CLIENTEMACTXDVLD ;
input CLIENTEMACTXDVLDMSW ;
input CLIENTEMACTXFIRSTBYTE ;
input CLIENTEMACTXUNDERRUN ;
input DCREMACCLK ;
input DCREMACENABLE ;
input DCREMACREAD ;
input DCREMACWRITE ;
input HOSTCLK ;
input HOSTMIIMSEL ;
input HOSTREQ ;
input PHYEMACCOL ;
input PHYEMACCRS ;
input PHYEMACGTXCLK ;
input PHYEMACMCLKIN ;
input PHYEMACMDIN ;
input PHYEMACMIITXCLK ;
input PHYEMACRXCHARISCOMMA ;
input PHYEMACRXCHARISK ;
input PHYEMACRXCLK ;
input PHYEMACRXDISPERR ;
input PHYEMACRXDV ;
input PHYEMACRXER ;
input PHYEMACRXNOTINTABLE ;
input PHYEMACRXRUNDISP ;
input PHYEMACSIGNALDET ;
input PHYEMACTXBUFERR ;
input PHYEMACTXGMIIMIICLKIN ;
input RESET ;
input [0:31] DCREMACDBUS ;
input [0:9] DCREMACABUS ;
input [15:0] CLIENTEMACPAUSEVAL ;
input [15:0] CLIENTEMACTXD ;
input [1:0] HOSTOPCODE ;
input [1:0] PHYEMACRXBUFSTATUS ;
input [2:0] PHYEMACRXCLKCORCNT ;
input [31:0] HOSTWRDATA ;
input [4:0] PHYEMACPHYAD ;
input [7:0] CLIENTEMACTXIFGDELAY ;
input [7:0] PHYEMACRXD ;
input [9:0] HOSTADDR ;
output DCRHOSTDONEIR ;
output EMACCLIENTANINTERRUPT ;
output EMACCLIENTRXBADFRAME ;
output EMACCLIENTRXCLIENTCLKOUT ;
output EMACCLIENTRXDVLD ;
output EMACCLIENTRXDVLDMSW ;
output EMACCLIENTRXFRAMEDROP ;
output EMACCLIENTRXGOODFRAME ;
output EMACCLIENTRXSTATSBYTEVLD ;
output EMACCLIENTRXSTATSVLD ;
output EMACCLIENTTXACK ;
output EMACCLIENTTXCLIENTCLKOUT ;
output EMACCLIENTTXCOLLISION ;
output EMACCLIENTTXRETRANSMIT ;
output EMACCLIENTTXSTATS ;
output EMACCLIENTTXSTATSBYTEVLD ;
output EMACCLIENTTXSTATSVLD ;
output EMACDCRACK ;
output EMACPHYENCOMMAALIGN ;
output EMACPHYLOOPBACKMSB ;
output EMACPHYMCLKOUT ;
output EMACPHYMDOUT ;
output EMACPHYMDTRI ;
output EMACPHYMGTRXRESET ;
output EMACPHYMGTTXRESET ;
output EMACPHYPOWERDOWN ;
output EMACPHYSYNCACQSTATUS ;
output EMACPHYTXCHARDISPMODE ;
output EMACPHYTXCHARDISPVAL ;
output EMACPHYTXCHARISK ;
output EMACPHYTXCLK ;
output EMACPHYTXEN ;
output EMACPHYTXER ;
output EMACPHYTXGMIIMIICLKOUT ;
output EMACSPEEDIS10100 ;
output HOSTMIIMRDY ;
output [0:31] EMACDCRDBUS ;
output [15:0] EMACCLIENTRXD ;
output [31:0] HOSTRDDATA ;
output [6:0] EMACCLIENTRXSTATS ;
output [7:0] EMACPHYTXD ;
parameter EMAC_1000BASEX_ENABLE = "FALSE";
parameter EMAC_ADDRFILTER_ENABLE = "FALSE";
parameter EMAC_BYTEPHY = "FALSE";
parameter EMAC_CTRLLENCHECK_DISABLE = "FALSE";
parameter [0:7] EMAC_DCRBASEADDR = 8'h00;
parameter EMAC_GTLOOPBACK = "FALSE";
parameter EMAC_HOST_ENABLE = "FALSE";
parameter [8:0] EMAC_LINKTIMERVAL = 9'h000;
parameter EMAC_LTCHECK_DISABLE = "FALSE";
parameter EMAC_MDIO_ENABLE = "FALSE";
parameter EMAC_MDIO_IGNORE_PHYADZERO = "FALSE";
parameter [47:0] EMAC_PAUSEADDR = 48'h000000000000;
parameter EMAC_PHYINITAUTONEG_ENABLE = "FALSE";
parameter EMAC_PHYISOLATE = "FALSE";
parameter EMAC_PHYLOOPBACKMSB = "FALSE";
parameter EMAC_PHYPOWERDOWN = "FALSE";
parameter EMAC_PHYRESET = "FALSE";
parameter EMAC_RGMII_ENABLE = "FALSE";
parameter EMAC_RX16BITCLIENT_ENABLE = "FALSE";
parameter EMAC_RXFLOWCTRL_ENABLE = "FALSE";
parameter EMAC_RXHALFDUPLEX = "FALSE";
parameter EMAC_RXINBANDFCS_ENABLE = "FALSE";
parameter EMAC_RXJUMBOFRAME_ENABLE = "FALSE";
parameter EMAC_RXRESET = "FALSE";
parameter EMAC_RXVLAN_ENABLE = "FALSE";
parameter EMAC_RX_ENABLE = "TRUE";
parameter EMAC_SGMII_ENABLE = "FALSE";
parameter EMAC_SPEED_LSB = "FALSE";
parameter EMAC_SPEED_MSB = "FALSE";
parameter EMAC_TX16BITCLIENT_ENABLE = "FALSE";
parameter EMAC_TXFLOWCTRL_ENABLE = "FALSE";
parameter EMAC_TXHALFDUPLEX = "FALSE";
parameter EMAC_TXIFGADJUST_ENABLE = "FALSE";
parameter EMAC_TXINBANDFCS_ENABLE = "FALSE";
parameter EMAC_TXJUMBOFRAME_ENABLE = "FALSE";
parameter EMAC_TXRESET = "FALSE";
parameter EMAC_TXVLAN_ENABLE = "FALSE";
parameter EMAC_TX_ENABLE = "TRUE";
parameter [47:0] EMAC_UNICASTADDR = 48'h000000000000;
parameter EMAC_UNIDIRECTION_ENABLE = "FALSE";
parameter EMAC_USECLKEN = "FALSE";
parameter SIM_VERSION = "1.0";
endmodule
//#### END MODULE DEFINITION FOR: TEMAC_SINGLE ####

//#### BEGIN MODULE DEFINITION FOR :TIMEGRP ###
module TIMEGRP () /* synthesis syn_black_box  syn_lib_cell=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: TIMEGRP ####

//#### BEGIN MODULE DEFINITION FOR :TIMESPEC ###
module TIMESPEC () /* synthesis syn_black_box  syn_lib_cell=1
 */;
endmodule
//#### END MODULE DEFINITION FOR: TIMESPEC ####

//#### BEGIN MODULE DEFINITION FOR :USR_ACCESSE2 ###
module USR_ACCESSE2 (
  CFGCLK,
  DATA,
  DATAVALID
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
output CFGCLK ;
output DATAVALID ;
output [31:0] DATA ;
endmodule
//#### END MODULE DEFINITION FOR: USR_ACCESSE2 ####

//#### BEGIN MODULE DEFINITION FOR :USR_ACCESS_VIRTEX4 ###
module USR_ACCESS_VIRTEX4 (DATA, DATAVALID) /* synthesis syn_black_box  syn_lib_cell=1
 */;
output [31:0] DATA ;
output DATAVALID ;
endmodule
//#### END MODULE DEFINITION FOR: USR_ACCESS_VIRTEX4 ####

//#### BEGIN MODULE DEFINITION FOR :USR_ACCESS_VIRTEX5 ###
module USR_ACCESS_VIRTEX5 (
        CFGCLK,
	DATA,
	DATAVALID
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
output CFGCLK ;
output DATAVALID ;
output [31:0] DATA ;
endmodule
//#### END MODULE DEFINITION FOR: USR_ACCESS_VIRTEX5 ####

//#### BEGIN MODULE DEFINITION FOR :USR_ACCESS_VIRTEX6 ###
module USR_ACCESS_VIRTEX6 (
  CFGCLK,
  DATA,
  DATAVALID
) /* synthesis syn_black_box  syn_lib_cell=1
 */;
output CFGCLK ;
output DATAVALID ;
output [31:0] DATA ;
endmodule
//#### END MODULE DEFINITION FOR: USR_ACCESS_VIRTEX6 ####

//#### BEGIN MODULE DEFINITION FOR :VCC ###
module VCC(P) /* synthesis syn_black_box  syn_lib_cell=1
 .noprune=1
 */;
output P ;
endmodule
//#### END MODULE DEFINITION FOR: VCC ####

//#### BEGIN MODULE DEFINITION FOR :XADC ###
module XADC (
        ALM,
        BUSY,
        CHANNEL,
        DO,
        DRDY,
        EOC,
        EOS,
        JTAGBUSY,
        JTAGLOCKED,
        JTAGMODIFIED,
        MUXADDR,
        OT,
        CONVST,
        CONVSTCLK,
        DADDR,
        DCLK,
        DEN,
        DI,
        DWE,
        RESET,
        VAUXN,
        VAUXP,
        VN,
        VP

) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CONVST ;
input CONVSTCLK ;
input DCLK ;
input DEN ;
input DWE ;
input RESET ;
input VN ;
input VP ;
input [15:0] DI ;
input [15:0] VAUXN ;
input [15:0] VAUXP ;
input [6:0] DADDR ;
output BUSY ;
output DRDY ;
output EOC ;
output EOS ;
output JTAGBUSY ;
output JTAGLOCKED ;
output JTAGMODIFIED ;
output OT ;
output [15:0] DO ;
output [7:0] ALM ;
output [4:0] CHANNEL ;
output [4:0] MUXADDR ;
parameter  [15:0] INIT_40 = 16'h0;
parameter  [15:0] INIT_41 = 16'h0;
parameter  [15:0] INIT_42 = 16'h0800;
parameter  [15:0] INIT_43 = 16'h0;
parameter  [15:0] INIT_44 = 16'h0;
parameter  [15:0] INIT_45 = 16'h0;
parameter  [15:0] INIT_46 = 16'h0;
parameter  [15:0] INIT_47 = 16'h0;
parameter  [15:0] INIT_48 = 16'h0;
parameter  [15:0] INIT_49 = 16'h0;
parameter  [15:0] INIT_4A = 16'h0;
parameter  [15:0] INIT_4B = 16'h0;
parameter  [15:0] INIT_4C = 16'h0;
parameter  [15:0] INIT_4D = 16'h0;
parameter  [15:0] INIT_4E = 16'h0;
parameter  [15:0] INIT_4F = 16'h0;
parameter  [15:0] INIT_50 = 16'h0;
parameter  [15:0] INIT_51 = 16'h0;
parameter  [15:0] INIT_52 = 16'h0;
parameter  [15:0] INIT_53 = 16'h0;
parameter  [15:0] INIT_54 = 16'h0;
parameter  [15:0] INIT_55 = 16'h0;
parameter  [15:0] INIT_56 = 16'h0;
parameter  [15:0] INIT_57 = 16'h0;
parameter  [15:0] INIT_58 = 16'h0;
parameter  [15:0] INIT_59 = 16'h0;
parameter  [15:0] INIT_5A = 16'h0;
parameter  [15:0] INIT_5B = 16'h0;
parameter  [15:0] INIT_5C = 16'h0;
parameter  [15:0] INIT_5D = 16'h0;
parameter  [15:0] INIT_5E = 16'h0;
parameter  [15:0] INIT_5F = 16'h0;
parameter SIM_DEVICE = "7SERIES";
parameter SIM_MONITOR_FILE = "design.txt";
endmodule
//#### END MODULE DEFINITION FOR: XADC ####

//#### BEGIN MODULE DEFINITION FOR :XNOR2 ###
module XNOR2 (O, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: XNOR2 ####

//#### BEGIN MODULE DEFINITION FOR :XNOR3 ###
module XNOR3 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: XNOR3 ####

//#### BEGIN MODULE DEFINITION FOR :XNOR4 ###
module XNOR4 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: XNOR4 ####

//#### BEGIN MODULE DEFINITION FOR :XNOR5 ###
module XNOR5 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: XNOR5 ####

//#### BEGIN MODULE DEFINITION FOR :XOR2 ###
module XOR2 (O, I0, I1) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: XOR2 ####

//#### BEGIN MODULE DEFINITION FOR :XOR3 ###
module XOR3 (O, I0, I1, I2) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: XOR3 ####

//#### BEGIN MODULE DEFINITION FOR :XOR4 ###
module XOR4 (O, I0, I1, I2, I3) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: XOR4 ####

//#### BEGIN MODULE DEFINITION FOR :XOR5 ###
module XOR5 (O, I0, I1, I2, I3, I4) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input I0 ;
input I1 ;
input I2 ;
input I3 ;
input I4 ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: XOR5 ####

//#### BEGIN MODULE DEFINITION FOR :XORCY ###
module XORCY (O, CI, LI) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CI ;
input LI ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: XORCY ####

//#### BEGIN MODULE DEFINITION FOR :XORCY_D ###
module XORCY_D (LO, O, CI, LI) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CI ;
input LI ;
output LO ;
output O ;
endmodule
//#### END MODULE DEFINITION FOR: XORCY_D ####

//#### BEGIN MODULE DEFINITION FOR :XORCY_L ###
module XORCY_L (LO, CI, LI) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input CI ;
input LI ;
output LO ;
endmodule
//#### END MODULE DEFINITION FOR: XORCY_L ####

//#### BEGIN MODULE DEFINITION FOR :ZHOLD_DELAY ###
module ZHOLD_DELAY (
          DLYFABRIC,
          DLYIFF,
          DLYIN
      ) /* synthesis syn_black_box  syn_lib_cell=1
 */;
input DLYIN ;
output DLYFABRIC ;
output DLYIFF ;
parameter ZHOLD_FABRIC = "DEFAULT";
parameter ZHOLD_IFF    = "DEFAULT";
endmodule
//#### END MODULE DEFINITION FOR: ZHOLD_DELAY ####

//####### Components added for backward compatibility #######
module IPAD (PAD) /* synthesis syn_black_box black_box_pad_pin = "PAD" */;
    output PAD;
endmodule

module OPAD (PAD) /* synthesis syn_black_box black_box_pad_pin = "PAD" */;
    input PAD;
endmodule
module STARTUP_VIRTEX2_CLK (CLK) /* synthesis syn_black_box .noprune=1 xc_alias="STARTUP_VIRTEX2"*/;
    input  CLK;
endmodule
module STARTUP_VIRTEX2_GSR (GSR) /* synthesis syn_black_box .noprune=1 xc_alias="STARTUP_VIRTEX2"*/;
    input  GSR;
endmodule
module STARTUP_VIRTEX2_GTS (GTS) /* synthesis syn_black_box .noprune=1 xc_alias="STARTUP_VIRTEX2"*/;
    input  GTS;
endmodule
module STARTUP_VIRTEX2_GHIGH (GHIGH) /* synthesis syn_black_box .noprune=1 xc_alias="STARTUP_VIRTEX2"*/;
    input  GHIGH;
endmodule
module STARTUP_VIRTEX2_GWE (GWE) /* synthesis syn_black_box .noprune=1 xc_alias="STARTUP_VIRTEX2"*/;
    input  GWE;
endmodule
module STARTUP_VIRTEX2_ALL(GSR, GTS, CLK)
/* synthesis syn_black_box .noprune=1 xc_alias="STARTUP_VIRTEX2" */ ;
input GSR /* synthesis syn_defaultvalue=0 */,
      GTS /* synthesis syn_defaultvalue=0 */,
      CLK /* synthesis syn_defaultvalue=0 */;
endmodule

module STARTUP_VIRTEX_CLK (CLK)
/* synthesis syn_black_box .noprune=1 xc_alias="STARTUP_VIRTEX"*/ ;
    input  CLK;
endmodule
module STARTUP_VIRTEX_GSR (GSR) /* synthesis syn_black_box .noprune=1 */;
    input  GSR;
endmodule
module STARTUP_VIRTEX_GTS (GTS) /* synthesis syn_black_box .noprune=1 xc_alias="STARTUP_VIRTEX"*/;
    input  GTS;
endmodule
module STARTUP_VIRTEX_ALL(GSR, GTS, CLK)
/* synthesis syn_black_box .noprune=1 xc_alias="STARTUP_VIRTEX" */ ;
input GSR /* synthesis syn_defaultvalue=0 */,
      GTS /* synthesis syn_defaultvalue=0 */,
      CLK /* synthesis syn_defaultvalue=0 */;
endmodule

module STARTUP_SPARTAN2_CLK (CLK)
/* synthesis syn_black_box .noprune=1 xc_alias="STARTUP_SPARTAN2"*/ ;
    input  CLK;
endmodule
module STARTUP_SPARTAN2_GSR (GSR) /* synthesis syn_black_box .noprune=1 */;
    input  GSR;
endmodule
module STARTUP_SPARTAN2_GTS (GTS) /* synthesis syn_black_box .noprune=1 xc_alias="STARTUP_SPARTAN2"*/;
    input  GTS;
endmodule
module STARTUP_SPARTAN2_ALL(GSR, GTS, CLK)
/* synthesis syn_black_box .noprune=1 xc_alias="STARTUP_SPARTAN2" */ ;
input GSR /* synthesis syn_defaultvalue=0 */,
      GTS /* synthesis syn_defaultvalue=0 */,
      CLK /* synthesis syn_defaultvalue=0 */;
endmodule
